module MMCME4_ADV_Wrapper(
  input   io_CLKIN1,
  output  io_LOCKED,
  output  io_CLKOUT0,
  output  io_CLKOUT1
);
  wire  mmcm4_adv_CLKIN1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKIN2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_RST; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PWRDWN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CDDCREQ; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKINSEL; // @[Buf.scala 109:25]
  wire [6:0] mmcm4_adv_DADDR; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DEN; // @[Buf.scala 109:25]
  wire [15:0] mmcm4_adv_DI; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DWE; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSEN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSINCDEC; // @[Buf.scala 109:25]
  wire  mmcm4_adv_LOCKED; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT0; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT3; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT4; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT5; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT6; // @[Buf.scala 109:25]
  MMCME4_ADV
    #(.CLKOUT5_DIVIDE(2), .CLKOUT3_DIVIDE(2), .CLKFBOUT_PHASE(0.0), .CLKIN1_PERIOD(10), .CLKOUT2_DIVIDE(12), .CLKOUT0_PHASE(0.0), .CLKFBOUT_MULT_F(12), .CLKOUT4_DIVIDE(2), .CLKOUT6_DIVIDE(2), .CLKOUT0_USE_FINE_PS("FALSE"), .COMPENSATION("INTERNAL"), .CLKOUT1_DIVIDE(4), .BANDWIDTH("OPTIMIZED"), .CLKFBOUT_USE_FINE_PS("FALSE"), .CLKOUT4_CASCADE("FALSE"), .CLKOUT0_DIVIDE_F(12), .CLKOUT0_DUTY_CYCLE(0.5), .REF_JITTER1(0.01), .DIVCLK_DIVIDE(1), .STARTUP_WAIT("FALSE"))
    mmcm4_adv ( // @[Buf.scala 109:25]
    .CLKIN1(mmcm4_adv_CLKIN1),
    .CLKIN2(mmcm4_adv_CLKIN2),
    .RST(mmcm4_adv_RST),
    .PWRDWN(mmcm4_adv_PWRDWN),
    .CDDCREQ(mmcm4_adv_CDDCREQ),
    .CLKINSEL(mmcm4_adv_CLKINSEL),
    .DADDR(mmcm4_adv_DADDR),
    .DEN(mmcm4_adv_DEN),
    .DI(mmcm4_adv_DI),
    .DWE(mmcm4_adv_DWE),
    .PSCLK(mmcm4_adv_PSCLK),
    .PSEN(mmcm4_adv_PSEN),
    .DCLK(mmcm4_adv_DCLK),
    .PSINCDEC(mmcm4_adv_PSINCDEC),
    .LOCKED(mmcm4_adv_LOCKED),
    .CLKOUT0(mmcm4_adv_CLKOUT0),
    .CLKOUT1(mmcm4_adv_CLKOUT1),
    .CLKOUT2(mmcm4_adv_CLKOUT2),
    .CLKOUT3(mmcm4_adv_CLKOUT3),
    .CLKOUT4(mmcm4_adv_CLKOUT4),
    .CLKOUT5(mmcm4_adv_CLKOUT5),
    .CLKOUT6(mmcm4_adv_CLKOUT6)
  );
  assign io_LOCKED = mmcm4_adv_LOCKED; // @[Buf.scala 123:26]
  assign io_CLKOUT0 = mmcm4_adv_CLKOUT0; // @[Buf.scala 124:26]
  assign io_CLKOUT1 = mmcm4_adv_CLKOUT1; // @[Buf.scala 125:26]
  assign mmcm4_adv_CLKIN1 = io_CLKIN1; // @[Buf.scala 121:26]
  assign mmcm4_adv_CLKIN2 = 1'h0; // @[Buf.scala 132:31]
  assign mmcm4_adv_RST = 1'h0; // @[Buf.scala 122:26]
  assign mmcm4_adv_PWRDWN = 1'h0; // @[Buf.scala 133:30]
  assign mmcm4_adv_CDDCREQ = 1'h0; // @[Buf.scala 134:32]
  assign mmcm4_adv_CLKINSEL = 1'h1; // @[Buf.scala 135:32]
  assign mmcm4_adv_DADDR = 7'h0; // @[Buf.scala 136:30]
  assign mmcm4_adv_DEN = 1'h0; // @[Buf.scala 137:28]
  assign mmcm4_adv_DI = 16'h0; // @[Buf.scala 138:26]
  assign mmcm4_adv_DWE = 1'h0; // @[Buf.scala 139:28]
  assign mmcm4_adv_PSCLK = 1'h0; // @[Buf.scala 140:30]
  assign mmcm4_adv_PSEN = 1'h0; // @[Buf.scala 141:28]
  assign mmcm4_adv_DCLK = 1'h0; // @[Buf.scala 142:28]
  assign mmcm4_adv_PSINCDEC = 1'h0; // @[Buf.scala 143:32]
endmodule
module MMCME4_ADV_Wrapper_1(
  input   io_CLKIN1,
  output  io_LOCKED,
  output  io_CLKOUT0,
  output  io_CLKOUT1,
  output  io_CLKOUT2,
  output  io_CLKOUT3,
  output  io_CLKOUT4,
  output  io_CLKOUT5
);
  wire  mmcm4_adv_CLKIN1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKIN2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_RST; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PWRDWN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CDDCREQ; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKINSEL; // @[Buf.scala 109:25]
  wire [6:0] mmcm4_adv_DADDR; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DEN; // @[Buf.scala 109:25]
  wire [15:0] mmcm4_adv_DI; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DWE; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSEN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSINCDEC; // @[Buf.scala 109:25]
  wire  mmcm4_adv_LOCKED; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT0; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT3; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT4; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT5; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT6; // @[Buf.scala 109:25]
  MMCME4_ADV
    #(.CLKOUT5_DIVIDE(12), .CLKOUT3_DIVIDE(12), .CLKFBOUT_PHASE(0.0), .CLKIN1_PERIOD(10), .CLKOUT2_DIVIDE(12), .CLKOUT0_PHASE(0.0), .CLKFBOUT_MULT_F(12), .CLKOUT4_DIVIDE(12), .CLKOUT6_DIVIDE(2), .CLKOUT0_USE_FINE_PS("FALSE"), .COMPENSATION("INTERNAL"), .CLKOUT1_DIVIDE(12), .BANDWIDTH("OPTIMIZED"), .CLKFBOUT_USE_FINE_PS("FALSE"), .CLKOUT4_CASCADE("FALSE"), .CLKOUT0_DIVIDE_F(12), .CLKOUT0_DUTY_CYCLE(0.5), .REF_JITTER1(0.01), .DIVCLK_DIVIDE(1), .STARTUP_WAIT("FALSE"))
    mmcm4_adv ( // @[Buf.scala 109:25]
    .CLKIN1(mmcm4_adv_CLKIN1),
    .CLKIN2(mmcm4_adv_CLKIN2),
    .RST(mmcm4_adv_RST),
    .PWRDWN(mmcm4_adv_PWRDWN),
    .CDDCREQ(mmcm4_adv_CDDCREQ),
    .CLKINSEL(mmcm4_adv_CLKINSEL),
    .DADDR(mmcm4_adv_DADDR),
    .DEN(mmcm4_adv_DEN),
    .DI(mmcm4_adv_DI),
    .DWE(mmcm4_adv_DWE),
    .PSCLK(mmcm4_adv_PSCLK),
    .PSEN(mmcm4_adv_PSEN),
    .DCLK(mmcm4_adv_DCLK),
    .PSINCDEC(mmcm4_adv_PSINCDEC),
    .LOCKED(mmcm4_adv_LOCKED),
    .CLKOUT0(mmcm4_adv_CLKOUT0),
    .CLKOUT1(mmcm4_adv_CLKOUT1),
    .CLKOUT2(mmcm4_adv_CLKOUT2),
    .CLKOUT3(mmcm4_adv_CLKOUT3),
    .CLKOUT4(mmcm4_adv_CLKOUT4),
    .CLKOUT5(mmcm4_adv_CLKOUT5),
    .CLKOUT6(mmcm4_adv_CLKOUT6)
  );
  assign io_LOCKED = mmcm4_adv_LOCKED; // @[Buf.scala 123:26]
  assign io_CLKOUT0 = mmcm4_adv_CLKOUT0; // @[Buf.scala 124:26]
  assign io_CLKOUT1 = mmcm4_adv_CLKOUT1; // @[Buf.scala 125:26]
  assign io_CLKOUT2 = mmcm4_adv_CLKOUT2; // @[Buf.scala 126:26]
  assign io_CLKOUT3 = mmcm4_adv_CLKOUT3; // @[Buf.scala 127:26]
  assign io_CLKOUT4 = mmcm4_adv_CLKOUT4; // @[Buf.scala 128:26]
  assign io_CLKOUT5 = mmcm4_adv_CLKOUT5; // @[Buf.scala 129:26]
  assign mmcm4_adv_CLKIN1 = io_CLKIN1; // @[Buf.scala 121:26]
  assign mmcm4_adv_CLKIN2 = 1'h0; // @[Buf.scala 132:31]
  assign mmcm4_adv_RST = 1'h0; // @[Buf.scala 122:26]
  assign mmcm4_adv_PWRDWN = 1'h0; // @[Buf.scala 133:30]
  assign mmcm4_adv_CDDCREQ = 1'h0; // @[Buf.scala 134:32]
  assign mmcm4_adv_CLKINSEL = 1'h1; // @[Buf.scala 135:32]
  assign mmcm4_adv_DADDR = 7'h0; // @[Buf.scala 136:30]
  assign mmcm4_adv_DEN = 1'h0; // @[Buf.scala 137:28]
  assign mmcm4_adv_DI = 16'h0; // @[Buf.scala 138:26]
  assign mmcm4_adv_DWE = 1'h0; // @[Buf.scala 139:28]
  assign mmcm4_adv_PSCLK = 1'h0; // @[Buf.scala 140:30]
  assign mmcm4_adv_PSEN = 1'h0; // @[Buf.scala 141:28]
  assign mmcm4_adv_DCLK = 1'h0; // @[Buf.scala 142:28]
  assign mmcm4_adv_PSINCDEC = 1'h0; // @[Buf.scala 143:32]
endmodule
module MMCME4_ADV_Wrapper_2(
  input   io_CLKIN1,
  input   io_RST,
  output  io_LOCKED,
  output  io_CLKOUT0
);
  wire  mmcm4_adv_CLKIN1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKIN2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_RST; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PWRDWN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CDDCREQ; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKINSEL; // @[Buf.scala 109:25]
  wire [6:0] mmcm4_adv_DADDR; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DEN; // @[Buf.scala 109:25]
  wire [15:0] mmcm4_adv_DI; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DWE; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSEN; // @[Buf.scala 109:25]
  wire  mmcm4_adv_DCLK; // @[Buf.scala 109:25]
  wire  mmcm4_adv_PSINCDEC; // @[Buf.scala 109:25]
  wire  mmcm4_adv_LOCKED; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT0; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT1; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT2; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT3; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT4; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT5; // @[Buf.scala 109:25]
  wire  mmcm4_adv_CLKOUT6; // @[Buf.scala 109:25]
  MMCME4_ADV
    #(.CLKOUT5_DIVIDE(2), .CLKOUT3_DIVIDE(2), .CLKFBOUT_PHASE(0.0), .CLKIN1_PERIOD(10), .CLKOUT2_DIVIDE(2), .CLKOUT0_PHASE(0.0), .CLKFBOUT_MULT_F(18), .CLKOUT4_DIVIDE(2), .CLKOUT6_DIVIDE(2), .CLKOUT0_USE_FINE_PS("FALSE"), .COMPENSATION("INTERNAL"), .CLKOUT1_DIVIDE(2), .BANDWIDTH("OPTIMIZED"), .CLKFBOUT_USE_FINE_PS("FALSE"), .CLKOUT4_CASCADE("FALSE"), .CLKOUT0_DIVIDE_F(2), .CLKOUT0_DUTY_CYCLE(0.5), .REF_JITTER1(0.01), .DIVCLK_DIVIDE(2), .STARTUP_WAIT("FALSE"))
    mmcm4_adv ( // @[Buf.scala 109:25]
    .CLKIN1(mmcm4_adv_CLKIN1),
    .CLKIN2(mmcm4_adv_CLKIN2),
    .RST(mmcm4_adv_RST),
    .PWRDWN(mmcm4_adv_PWRDWN),
    .CDDCREQ(mmcm4_adv_CDDCREQ),
    .CLKINSEL(mmcm4_adv_CLKINSEL),
    .DADDR(mmcm4_adv_DADDR),
    .DEN(mmcm4_adv_DEN),
    .DI(mmcm4_adv_DI),
    .DWE(mmcm4_adv_DWE),
    .PSCLK(mmcm4_adv_PSCLK),
    .PSEN(mmcm4_adv_PSEN),
    .DCLK(mmcm4_adv_DCLK),
    .PSINCDEC(mmcm4_adv_PSINCDEC),
    .LOCKED(mmcm4_adv_LOCKED),
    .CLKOUT0(mmcm4_adv_CLKOUT0),
    .CLKOUT1(mmcm4_adv_CLKOUT1),
    .CLKOUT2(mmcm4_adv_CLKOUT2),
    .CLKOUT3(mmcm4_adv_CLKOUT3),
    .CLKOUT4(mmcm4_adv_CLKOUT4),
    .CLKOUT5(mmcm4_adv_CLKOUT5),
    .CLKOUT6(mmcm4_adv_CLKOUT6)
  );
  assign io_LOCKED = mmcm4_adv_LOCKED; // @[Buf.scala 123:26]
  assign io_CLKOUT0 = mmcm4_adv_CLKOUT0; // @[Buf.scala 124:26]
  assign mmcm4_adv_CLKIN1 = io_CLKIN1; // @[Buf.scala 121:26]
  assign mmcm4_adv_CLKIN2 = 1'h0; // @[Buf.scala 132:31]
  assign mmcm4_adv_RST = io_RST; // @[Buf.scala 122:26]
  assign mmcm4_adv_PWRDWN = 1'h0; // @[Buf.scala 133:30]
  assign mmcm4_adv_CDDCREQ = 1'h0; // @[Buf.scala 134:32]
  assign mmcm4_adv_CLKINSEL = 1'h1; // @[Buf.scala 135:32]
  assign mmcm4_adv_DADDR = 7'h0; // @[Buf.scala 136:30]
  assign mmcm4_adv_DEN = 1'h0; // @[Buf.scala 137:28]
  assign mmcm4_adv_DI = 16'h0; // @[Buf.scala 138:26]
  assign mmcm4_adv_DWE = 1'h0; // @[Buf.scala 139:28]
  assign mmcm4_adv_PSCLK = 1'h0; // @[Buf.scala 140:30]
  assign mmcm4_adv_PSEN = 1'h0; // @[Buf.scala 141:28]
  assign mmcm4_adv_DCLK = 1'h0; // @[Buf.scala 142:28]
  assign mmcm4_adv_PSINCDEC = 1'h0; // @[Buf.scala 143:32]
endmodule
module HBM_DRIVER(
  input          clock,
  output         io_hbm_clk,
  output         io_hbm_rstn,
  output         io_axi_hbm_0_aw_ready,
  input          io_axi_hbm_0_aw_valid,
  input  [33:0]  io_axi_hbm_0_aw_bits_addr,
  input  [3:0]   io_axi_hbm_0_aw_bits_len,
  output         io_axi_hbm_0_ar_ready,
  input          io_axi_hbm_0_ar_valid,
  input  [33:0]  io_axi_hbm_0_ar_bits_addr,
  input  [3:0]   io_axi_hbm_0_ar_bits_len,
  output         io_axi_hbm_0_w_ready,
  input          io_axi_hbm_0_w_valid,
  input  [255:0] io_axi_hbm_0_w_bits_data,
  input          io_axi_hbm_0_w_bits_last,
  input          io_axi_hbm_0_r_ready,
  output         io_axi_hbm_0_r_valid,
  output [255:0] io_axi_hbm_0_r_bits_data,
  output         io_axi_hbm_1_aw_ready,
  input          io_axi_hbm_1_aw_valid,
  input  [33:0]  io_axi_hbm_1_aw_bits_addr,
  input  [1:0]   io_axi_hbm_1_aw_bits_burst,
  input  [3:0]   io_axi_hbm_1_aw_bits_len,
  input  [2:0]   io_axi_hbm_1_aw_bits_size,
  output         io_axi_hbm_1_ar_ready,
  input          io_axi_hbm_1_ar_valid,
  input  [33:0]  io_axi_hbm_1_ar_bits_addr,
  input  [1:0]   io_axi_hbm_1_ar_bits_burst,
  input  [3:0]   io_axi_hbm_1_ar_bits_len,
  input  [2:0]   io_axi_hbm_1_ar_bits_size,
  output         io_axi_hbm_1_w_ready,
  input          io_axi_hbm_1_w_valid,
  input  [255:0] io_axi_hbm_1_w_bits_data,
  input          io_axi_hbm_1_w_bits_last,
  input  [31:0]  io_axi_hbm_1_w_bits_strb,
  input          io_axi_hbm_1_r_ready,
  output         io_axi_hbm_1_r_valid,
  output [255:0] io_axi_hbm_1_r_bits_data,
  output         io_axi_hbm_1_r_bits_last,
  input          io_axi_hbm_1_b_ready,
  output         io_axi_hbm_1_b_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  mmcmGlbl_io_CLKIN1; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_LOCKED; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT0; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT1; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT2; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT3; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT4; // @[HBMDriver.scala 48:30]
  wire  mmcmGlbl_io_CLKOUT5; // @[HBMDriver.scala 48:30]
  wire  apb0Pclk_pad_O; // @[Buf.scala 33:34]
  wire  apb0Pclk_pad_I; // @[Buf.scala 33:34]
  wire  apb0Pclk_pad_1_O; // @[Buf.scala 17:34]
  wire  apb0Pclk_pad_1_I; // @[Buf.scala 17:34]
  wire  apb0Pclk_pad_2_O; // @[Buf.scala 33:34]
  wire  apb0Pclk_pad_2_I; // @[Buf.scala 33:34]
  wire  axiAclkIn0_pad_O; // @[Buf.scala 33:34]
  wire  axiAclkIn0_pad_I; // @[Buf.scala 33:34]
  wire  hbmRefClk0_pad_O; // @[Buf.scala 33:34]
  wire  hbmRefClk0_pad_I; // @[Buf.scala 33:34]
  wire  apb1Pclk_pad_O; // @[Buf.scala 33:34]
  wire  apb1Pclk_pad_I; // @[Buf.scala 33:34]
  wire  apb1Pclk_pad_1_O; // @[Buf.scala 17:34]
  wire  apb1Pclk_pad_1_I; // @[Buf.scala 17:34]
  wire  apb1Pclk_pad_2_O; // @[Buf.scala 33:34]
  wire  apb1Pclk_pad_2_I; // @[Buf.scala 33:34]
  wire  axiAclkIn1_pad_O; // @[Buf.scala 33:34]
  wire  axiAclkIn1_pad_I; // @[Buf.scala 33:34]
  wire  hbmRefClk1_pad_O; // @[Buf.scala 33:34]
  wire  hbmRefClk1_pad_I; // @[Buf.scala 33:34]
  wire  mmcmAxi_io_CLKIN1; // @[HBMDriver.scala 71:29]
  wire  mmcmAxi_io_RST; // @[HBMDriver.scala 71:29]
  wire  mmcmAxi_io_LOCKED; // @[HBMDriver.scala 71:29]
  wire  mmcmAxi_io_CLKOUT0; // @[HBMDriver.scala 71:29]
  wire  axiAclk_pad_O; // @[Buf.scala 33:34]
  wire  axiAclk_pad_I; // @[Buf.scala 33:34]
  wire  instHbm_HBM_REF_CLK_0; // @[HBMDriver.scala 92:29]
  wire  instHbm_HBM_REF_CLK_1; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_00_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_00_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_00_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_00_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_00_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_00_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_00_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_00_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_00_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_00_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_00_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_00_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_00_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_00_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_00_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_00_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_00_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_00_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_00_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_00_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_01_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_01_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_01_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_01_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_01_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_01_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_01_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_01_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_01_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_01_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_01_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_01_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_01_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_01_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_01_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_01_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_01_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_01_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_01_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_01_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_02_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_02_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_02_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_02_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_02_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_02_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_02_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_02_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_02_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_02_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_02_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_02_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_02_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_02_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_02_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_02_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_02_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_02_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_02_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_02_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_03_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_03_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_03_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_03_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_03_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_03_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_03_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_03_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_03_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_03_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_03_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_03_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_03_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_03_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_03_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_03_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_03_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_03_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_03_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_03_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_04_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_04_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_04_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_04_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_04_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_04_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_04_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_04_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_04_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_04_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_04_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_04_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_04_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_04_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_04_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_04_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_04_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_04_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_04_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_04_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_05_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_05_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_05_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_05_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_05_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_05_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_05_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_05_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_05_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_05_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_05_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_05_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_05_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_05_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_05_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_05_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_05_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_05_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_05_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_05_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_06_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_06_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_06_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_06_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_06_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_06_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_06_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_06_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_06_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_06_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_06_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_06_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_06_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_06_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_06_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_06_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_06_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_06_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_06_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_06_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_07_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_07_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_07_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_07_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_07_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_07_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_07_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_07_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_07_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_07_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_07_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_07_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_07_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_07_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_07_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_07_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_07_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_07_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_07_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_07_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_08_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_08_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_08_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_08_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_08_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_08_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_08_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_08_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_08_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_08_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_08_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_08_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_08_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_08_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_08_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_08_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_08_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_08_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_08_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_08_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_09_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_09_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_09_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_09_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_09_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_09_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_09_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_09_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_09_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_09_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_09_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_09_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_09_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_09_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_09_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_09_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_09_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_09_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_09_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_09_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_10_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_10_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_10_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_10_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_10_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_10_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_10_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_10_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_10_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_10_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_10_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_10_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_10_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_10_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_10_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_10_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_10_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_10_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_10_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_10_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_11_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_11_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_11_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_11_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_11_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_11_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_11_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_11_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_11_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_11_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_11_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_11_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_11_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_11_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_11_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_11_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_11_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_11_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_11_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_11_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_12_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_12_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_12_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_12_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_12_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_12_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_12_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_12_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_12_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_12_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_12_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_12_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_12_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_12_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_12_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_12_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_12_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_12_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_12_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_12_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_13_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_13_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_13_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_13_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_13_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_13_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_13_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_13_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_13_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_13_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_13_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_13_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_13_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_13_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_13_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_13_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_13_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_13_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_13_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_13_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_14_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_14_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_14_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_14_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_14_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_14_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_14_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_14_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_14_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_14_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_14_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_14_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_14_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_14_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_14_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_14_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_14_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_14_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_14_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_14_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_15_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_15_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_15_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_15_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_15_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_15_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_15_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_15_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_15_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_15_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_15_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_15_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_15_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_15_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_15_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_15_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_15_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_15_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_15_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_15_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_16_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_16_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_16_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_16_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_16_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_16_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_16_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_16_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_16_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_16_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_16_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_16_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_16_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_16_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_16_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_16_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_16_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_16_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_16_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_16_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_17_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_17_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_17_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_17_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_17_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_17_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_17_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_17_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_17_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_17_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_17_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_17_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_17_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_17_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_17_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_17_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_17_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_17_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_17_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_17_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_18_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_18_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_18_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_18_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_18_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_18_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_18_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_18_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_18_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_18_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_18_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_18_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_18_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_18_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_18_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_18_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_18_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_18_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_18_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_18_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_19_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_19_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_19_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_19_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_19_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_19_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_19_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_19_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_19_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_19_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_19_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_19_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_19_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_19_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_19_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_19_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_19_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_19_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_19_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_19_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_20_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_20_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_20_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_20_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_20_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_20_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_20_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_20_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_20_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_20_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_20_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_20_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_20_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_20_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_20_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_20_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_20_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_20_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_20_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_20_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_21_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_21_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_21_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_21_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_21_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_21_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_21_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_21_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_21_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_21_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_21_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_21_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_21_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_21_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_21_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_21_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_21_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_21_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_21_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_21_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_22_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_22_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_22_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_22_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_22_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_22_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_22_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_22_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_22_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_22_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_22_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_22_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_22_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_22_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_22_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_22_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_22_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_22_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_22_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_22_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_23_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_23_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_23_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_23_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_23_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_23_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_23_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_23_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_23_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_23_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_23_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_23_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_23_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_23_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_23_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_23_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_23_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_23_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_23_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_23_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_24_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_24_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_24_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_24_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_24_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_24_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_24_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_24_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_24_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_24_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_24_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_24_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_24_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_24_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_24_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_24_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_24_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_24_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_24_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_24_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_25_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_25_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_25_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_25_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_25_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_25_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_25_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_25_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_25_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_25_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_25_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_25_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_25_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_25_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_25_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_25_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_25_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_25_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_25_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_25_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_26_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_26_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_26_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_26_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_26_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_26_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_26_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_26_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_26_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_26_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_26_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_26_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_26_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_26_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_26_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_26_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_26_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_26_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_26_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_26_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_27_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_27_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_27_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_27_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_27_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_27_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_27_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_27_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_27_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_27_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_27_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_27_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_27_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_27_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_27_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_27_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_27_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_27_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_27_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_27_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_28_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_28_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_28_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_28_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_28_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_28_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_28_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_28_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_28_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_28_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_28_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_28_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_28_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_28_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_28_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_28_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_28_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_28_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_28_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_28_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_29_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_29_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_29_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_29_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_29_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_29_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_29_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_29_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_29_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_29_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_29_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_29_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_29_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_29_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_29_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_29_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_29_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_29_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_29_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_29_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_30_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_30_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_30_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_30_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_30_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_30_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_30_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_30_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_30_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_30_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_30_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_30_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_30_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_30_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_30_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_30_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_30_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_30_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_30_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_30_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_ACLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_ARESET_N; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_31_ARADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_31_ARBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_31_ARID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_31_ARLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_31_ARSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_ARVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_ARREADY; // @[HBMDriver.scala 92:29]
  wire [32:0] instHbm_AXI_31_AWADDR; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_31_AWBURST; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_31_AWID; // @[HBMDriver.scala 92:29]
  wire [3:0] instHbm_AXI_31_AWLEN; // @[HBMDriver.scala 92:29]
  wire [2:0] instHbm_AXI_31_AWSIZE; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_AWVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_AWREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_31_WDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_WLAST; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_31_WSTRB; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_WVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_WREADY; // @[HBMDriver.scala 92:29]
  wire [255:0] instHbm_AXI_31_RDATA; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_31_RID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_RLAST; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_31_RRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_RVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_RREADY; // @[HBMDriver.scala 92:29]
  wire [5:0] instHbm_AXI_31_BID; // @[HBMDriver.scala 92:29]
  wire [1:0] instHbm_AXI_31_BRESP; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_BVALID; // @[HBMDriver.scala 92:29]
  wire  instHbm_AXI_31_BREADY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_31_WDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_AXI_31_RDATA_PARITY; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_APB_0_PWDATA; // @[HBMDriver.scala 92:29]
  wire [21:0] instHbm_APB_0_PADDR; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PCLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PENABLE; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PRESET_N; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PSEL; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PWRITE; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_APB_0_PRDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PREADY; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_0_PSLVERR; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_APB_1_PWDATA; // @[HBMDriver.scala 92:29]
  wire [21:0] instHbm_APB_1_PADDR; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PCLK; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PENABLE; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PRESET_N; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PSEL; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PWRITE; // @[HBMDriver.scala 92:29]
  wire [31:0] instHbm_APB_1_PRDATA; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PREADY; // @[HBMDriver.scala 92:29]
  wire  instHbm_APB_1_PSLVERR; // @[HBMDriver.scala 92:29]
  wire  instHbm_DRAM_0_STAT_CATTRIP; // @[HBMDriver.scala 92:29]
  wire [6:0] instHbm_DRAM_0_STAT_TEMP; // @[HBMDriver.scala 92:29]
  wire  instHbm_DRAM_1_STAT_CATTRIP; // @[HBMDriver.scala 92:29]
  wire [6:0] instHbm_DRAM_1_STAT_TEMP; // @[HBMDriver.scala 92:29]
  wire  instHbm_apb_complete_0; // @[HBMDriver.scala 92:29]
  wire  instHbm_apb_complete_1; // @[HBMDriver.scala 92:29]
  reg  apb_complete_0_r; // @[Reg.scala 15:16]
  reg  apb_complete_0; // @[Reg.scala 15:16]
  reg  apb_complete_1_r; // @[Reg.scala 15:16]
  reg  apb_complete_1; // @[Reg.scala 15:16]
  reg  io_hbm_rstn_REG; // @[HBMDriver.scala 97:52]
  wire  _io_hbm_rstn_T_2 = io_hbm_rstn_REG & apb_complete_0; // @[HBMDriver.scala 98:17]
  MMCME4_ADV_Wrapper_1 mmcmGlbl ( // @[HBMDriver.scala 48:30]
    .io_CLKIN1(mmcmGlbl_io_CLKIN1),
    .io_LOCKED(mmcmGlbl_io_LOCKED),
    .io_CLKOUT0(mmcmGlbl_io_CLKOUT0),
    .io_CLKOUT1(mmcmGlbl_io_CLKOUT1),
    .io_CLKOUT2(mmcmGlbl_io_CLKOUT2),
    .io_CLKOUT3(mmcmGlbl_io_CLKOUT3),
    .io_CLKOUT4(mmcmGlbl_io_CLKOUT4),
    .io_CLKOUT5(mmcmGlbl_io_CLKOUT5)
  );
  BUFG apb0Pclk_pad ( // @[Buf.scala 33:34]
    .O(apb0Pclk_pad_O),
    .I(apb0Pclk_pad_I)
  );
  IBUF apb0Pclk_pad_1 ( // @[Buf.scala 17:34]
    .O(apb0Pclk_pad_1_O),
    .I(apb0Pclk_pad_1_I)
  );
  BUFG apb0Pclk_pad_2 ( // @[Buf.scala 33:34]
    .O(apb0Pclk_pad_2_O),
    .I(apb0Pclk_pad_2_I)
  );
  BUFG axiAclkIn0_pad ( // @[Buf.scala 33:34]
    .O(axiAclkIn0_pad_O),
    .I(axiAclkIn0_pad_I)
  );
  BUFG hbmRefClk0_pad ( // @[Buf.scala 33:34]
    .O(hbmRefClk0_pad_O),
    .I(hbmRefClk0_pad_I)
  );
  BUFG apb1Pclk_pad ( // @[Buf.scala 33:34]
    .O(apb1Pclk_pad_O),
    .I(apb1Pclk_pad_I)
  );
  IBUF apb1Pclk_pad_1 ( // @[Buf.scala 17:34]
    .O(apb1Pclk_pad_1_O),
    .I(apb1Pclk_pad_1_I)
  );
  BUFG apb1Pclk_pad_2 ( // @[Buf.scala 33:34]
    .O(apb1Pclk_pad_2_O),
    .I(apb1Pclk_pad_2_I)
  );
  BUFG axiAclkIn1_pad ( // @[Buf.scala 33:34]
    .O(axiAclkIn1_pad_O),
    .I(axiAclkIn1_pad_I)
  );
  BUFG hbmRefClk1_pad ( // @[Buf.scala 33:34]
    .O(hbmRefClk1_pad_O),
    .I(hbmRefClk1_pad_I)
  );
  MMCME4_ADV_Wrapper_2 mmcmAxi ( // @[HBMDriver.scala 71:29]
    .io_CLKIN1(mmcmAxi_io_CLKIN1),
    .io_RST(mmcmAxi_io_RST),
    .io_LOCKED(mmcmAxi_io_LOCKED),
    .io_CLKOUT0(mmcmAxi_io_CLKOUT0)
  );
  BUFG axiAclk_pad ( // @[Buf.scala 33:34]
    .O(axiAclk_pad_O),
    .I(axiAclk_pad_I)
  );
  HBMBlackBox instHbm ( // @[HBMDriver.scala 92:29]
    .HBM_REF_CLK_0(instHbm_HBM_REF_CLK_0),
    .HBM_REF_CLK_1(instHbm_HBM_REF_CLK_1),
    .AXI_00_ACLK(instHbm_AXI_00_ACLK),
    .AXI_00_ARESET_N(instHbm_AXI_00_ARESET_N),
    .AXI_00_ARADDR(instHbm_AXI_00_ARADDR),
    .AXI_00_ARBURST(instHbm_AXI_00_ARBURST),
    .AXI_00_ARID(instHbm_AXI_00_ARID),
    .AXI_00_ARLEN(instHbm_AXI_00_ARLEN),
    .AXI_00_ARSIZE(instHbm_AXI_00_ARSIZE),
    .AXI_00_ARVALID(instHbm_AXI_00_ARVALID),
    .AXI_00_ARREADY(instHbm_AXI_00_ARREADY),
    .AXI_00_AWADDR(instHbm_AXI_00_AWADDR),
    .AXI_00_AWBURST(instHbm_AXI_00_AWBURST),
    .AXI_00_AWID(instHbm_AXI_00_AWID),
    .AXI_00_AWLEN(instHbm_AXI_00_AWLEN),
    .AXI_00_AWSIZE(instHbm_AXI_00_AWSIZE),
    .AXI_00_AWVALID(instHbm_AXI_00_AWVALID),
    .AXI_00_AWREADY(instHbm_AXI_00_AWREADY),
    .AXI_00_WDATA(instHbm_AXI_00_WDATA),
    .AXI_00_WLAST(instHbm_AXI_00_WLAST),
    .AXI_00_WSTRB(instHbm_AXI_00_WSTRB),
    .AXI_00_WVALID(instHbm_AXI_00_WVALID),
    .AXI_00_WREADY(instHbm_AXI_00_WREADY),
    .AXI_00_RDATA(instHbm_AXI_00_RDATA),
    .AXI_00_RID(instHbm_AXI_00_RID),
    .AXI_00_RLAST(instHbm_AXI_00_RLAST),
    .AXI_00_RRESP(instHbm_AXI_00_RRESP),
    .AXI_00_RVALID(instHbm_AXI_00_RVALID),
    .AXI_00_RREADY(instHbm_AXI_00_RREADY),
    .AXI_00_BID(instHbm_AXI_00_BID),
    .AXI_00_BRESP(instHbm_AXI_00_BRESP),
    .AXI_00_BVALID(instHbm_AXI_00_BVALID),
    .AXI_00_BREADY(instHbm_AXI_00_BREADY),
    .AXI_00_WDATA_PARITY(instHbm_AXI_00_WDATA_PARITY),
    .AXI_00_RDATA_PARITY(instHbm_AXI_00_RDATA_PARITY),
    .AXI_01_ACLK(instHbm_AXI_01_ACLK),
    .AXI_01_ARESET_N(instHbm_AXI_01_ARESET_N),
    .AXI_01_ARADDR(instHbm_AXI_01_ARADDR),
    .AXI_01_ARBURST(instHbm_AXI_01_ARBURST),
    .AXI_01_ARID(instHbm_AXI_01_ARID),
    .AXI_01_ARLEN(instHbm_AXI_01_ARLEN),
    .AXI_01_ARSIZE(instHbm_AXI_01_ARSIZE),
    .AXI_01_ARVALID(instHbm_AXI_01_ARVALID),
    .AXI_01_ARREADY(instHbm_AXI_01_ARREADY),
    .AXI_01_AWADDR(instHbm_AXI_01_AWADDR),
    .AXI_01_AWBURST(instHbm_AXI_01_AWBURST),
    .AXI_01_AWID(instHbm_AXI_01_AWID),
    .AXI_01_AWLEN(instHbm_AXI_01_AWLEN),
    .AXI_01_AWSIZE(instHbm_AXI_01_AWSIZE),
    .AXI_01_AWVALID(instHbm_AXI_01_AWVALID),
    .AXI_01_AWREADY(instHbm_AXI_01_AWREADY),
    .AXI_01_WDATA(instHbm_AXI_01_WDATA),
    .AXI_01_WLAST(instHbm_AXI_01_WLAST),
    .AXI_01_WSTRB(instHbm_AXI_01_WSTRB),
    .AXI_01_WVALID(instHbm_AXI_01_WVALID),
    .AXI_01_WREADY(instHbm_AXI_01_WREADY),
    .AXI_01_RDATA(instHbm_AXI_01_RDATA),
    .AXI_01_RID(instHbm_AXI_01_RID),
    .AXI_01_RLAST(instHbm_AXI_01_RLAST),
    .AXI_01_RRESP(instHbm_AXI_01_RRESP),
    .AXI_01_RVALID(instHbm_AXI_01_RVALID),
    .AXI_01_RREADY(instHbm_AXI_01_RREADY),
    .AXI_01_BID(instHbm_AXI_01_BID),
    .AXI_01_BRESP(instHbm_AXI_01_BRESP),
    .AXI_01_BVALID(instHbm_AXI_01_BVALID),
    .AXI_01_BREADY(instHbm_AXI_01_BREADY),
    .AXI_01_WDATA_PARITY(instHbm_AXI_01_WDATA_PARITY),
    .AXI_01_RDATA_PARITY(instHbm_AXI_01_RDATA_PARITY),
    .AXI_02_ACLK(instHbm_AXI_02_ACLK),
    .AXI_02_ARESET_N(instHbm_AXI_02_ARESET_N),
    .AXI_02_ARADDR(instHbm_AXI_02_ARADDR),
    .AXI_02_ARBURST(instHbm_AXI_02_ARBURST),
    .AXI_02_ARID(instHbm_AXI_02_ARID),
    .AXI_02_ARLEN(instHbm_AXI_02_ARLEN),
    .AXI_02_ARSIZE(instHbm_AXI_02_ARSIZE),
    .AXI_02_ARVALID(instHbm_AXI_02_ARVALID),
    .AXI_02_ARREADY(instHbm_AXI_02_ARREADY),
    .AXI_02_AWADDR(instHbm_AXI_02_AWADDR),
    .AXI_02_AWBURST(instHbm_AXI_02_AWBURST),
    .AXI_02_AWID(instHbm_AXI_02_AWID),
    .AXI_02_AWLEN(instHbm_AXI_02_AWLEN),
    .AXI_02_AWSIZE(instHbm_AXI_02_AWSIZE),
    .AXI_02_AWVALID(instHbm_AXI_02_AWVALID),
    .AXI_02_AWREADY(instHbm_AXI_02_AWREADY),
    .AXI_02_WDATA(instHbm_AXI_02_WDATA),
    .AXI_02_WLAST(instHbm_AXI_02_WLAST),
    .AXI_02_WSTRB(instHbm_AXI_02_WSTRB),
    .AXI_02_WVALID(instHbm_AXI_02_WVALID),
    .AXI_02_WREADY(instHbm_AXI_02_WREADY),
    .AXI_02_RDATA(instHbm_AXI_02_RDATA),
    .AXI_02_RID(instHbm_AXI_02_RID),
    .AXI_02_RLAST(instHbm_AXI_02_RLAST),
    .AXI_02_RRESP(instHbm_AXI_02_RRESP),
    .AXI_02_RVALID(instHbm_AXI_02_RVALID),
    .AXI_02_RREADY(instHbm_AXI_02_RREADY),
    .AXI_02_BID(instHbm_AXI_02_BID),
    .AXI_02_BRESP(instHbm_AXI_02_BRESP),
    .AXI_02_BVALID(instHbm_AXI_02_BVALID),
    .AXI_02_BREADY(instHbm_AXI_02_BREADY),
    .AXI_02_WDATA_PARITY(instHbm_AXI_02_WDATA_PARITY),
    .AXI_02_RDATA_PARITY(instHbm_AXI_02_RDATA_PARITY),
    .AXI_03_ACLK(instHbm_AXI_03_ACLK),
    .AXI_03_ARESET_N(instHbm_AXI_03_ARESET_N),
    .AXI_03_ARADDR(instHbm_AXI_03_ARADDR),
    .AXI_03_ARBURST(instHbm_AXI_03_ARBURST),
    .AXI_03_ARID(instHbm_AXI_03_ARID),
    .AXI_03_ARLEN(instHbm_AXI_03_ARLEN),
    .AXI_03_ARSIZE(instHbm_AXI_03_ARSIZE),
    .AXI_03_ARVALID(instHbm_AXI_03_ARVALID),
    .AXI_03_ARREADY(instHbm_AXI_03_ARREADY),
    .AXI_03_AWADDR(instHbm_AXI_03_AWADDR),
    .AXI_03_AWBURST(instHbm_AXI_03_AWBURST),
    .AXI_03_AWID(instHbm_AXI_03_AWID),
    .AXI_03_AWLEN(instHbm_AXI_03_AWLEN),
    .AXI_03_AWSIZE(instHbm_AXI_03_AWSIZE),
    .AXI_03_AWVALID(instHbm_AXI_03_AWVALID),
    .AXI_03_AWREADY(instHbm_AXI_03_AWREADY),
    .AXI_03_WDATA(instHbm_AXI_03_WDATA),
    .AXI_03_WLAST(instHbm_AXI_03_WLAST),
    .AXI_03_WSTRB(instHbm_AXI_03_WSTRB),
    .AXI_03_WVALID(instHbm_AXI_03_WVALID),
    .AXI_03_WREADY(instHbm_AXI_03_WREADY),
    .AXI_03_RDATA(instHbm_AXI_03_RDATA),
    .AXI_03_RID(instHbm_AXI_03_RID),
    .AXI_03_RLAST(instHbm_AXI_03_RLAST),
    .AXI_03_RRESP(instHbm_AXI_03_RRESP),
    .AXI_03_RVALID(instHbm_AXI_03_RVALID),
    .AXI_03_RREADY(instHbm_AXI_03_RREADY),
    .AXI_03_BID(instHbm_AXI_03_BID),
    .AXI_03_BRESP(instHbm_AXI_03_BRESP),
    .AXI_03_BVALID(instHbm_AXI_03_BVALID),
    .AXI_03_BREADY(instHbm_AXI_03_BREADY),
    .AXI_03_WDATA_PARITY(instHbm_AXI_03_WDATA_PARITY),
    .AXI_03_RDATA_PARITY(instHbm_AXI_03_RDATA_PARITY),
    .AXI_04_ACLK(instHbm_AXI_04_ACLK),
    .AXI_04_ARESET_N(instHbm_AXI_04_ARESET_N),
    .AXI_04_ARADDR(instHbm_AXI_04_ARADDR),
    .AXI_04_ARBURST(instHbm_AXI_04_ARBURST),
    .AXI_04_ARID(instHbm_AXI_04_ARID),
    .AXI_04_ARLEN(instHbm_AXI_04_ARLEN),
    .AXI_04_ARSIZE(instHbm_AXI_04_ARSIZE),
    .AXI_04_ARVALID(instHbm_AXI_04_ARVALID),
    .AXI_04_ARREADY(instHbm_AXI_04_ARREADY),
    .AXI_04_AWADDR(instHbm_AXI_04_AWADDR),
    .AXI_04_AWBURST(instHbm_AXI_04_AWBURST),
    .AXI_04_AWID(instHbm_AXI_04_AWID),
    .AXI_04_AWLEN(instHbm_AXI_04_AWLEN),
    .AXI_04_AWSIZE(instHbm_AXI_04_AWSIZE),
    .AXI_04_AWVALID(instHbm_AXI_04_AWVALID),
    .AXI_04_AWREADY(instHbm_AXI_04_AWREADY),
    .AXI_04_WDATA(instHbm_AXI_04_WDATA),
    .AXI_04_WLAST(instHbm_AXI_04_WLAST),
    .AXI_04_WSTRB(instHbm_AXI_04_WSTRB),
    .AXI_04_WVALID(instHbm_AXI_04_WVALID),
    .AXI_04_WREADY(instHbm_AXI_04_WREADY),
    .AXI_04_RDATA(instHbm_AXI_04_RDATA),
    .AXI_04_RID(instHbm_AXI_04_RID),
    .AXI_04_RLAST(instHbm_AXI_04_RLAST),
    .AXI_04_RRESP(instHbm_AXI_04_RRESP),
    .AXI_04_RVALID(instHbm_AXI_04_RVALID),
    .AXI_04_RREADY(instHbm_AXI_04_RREADY),
    .AXI_04_BID(instHbm_AXI_04_BID),
    .AXI_04_BRESP(instHbm_AXI_04_BRESP),
    .AXI_04_BVALID(instHbm_AXI_04_BVALID),
    .AXI_04_BREADY(instHbm_AXI_04_BREADY),
    .AXI_04_WDATA_PARITY(instHbm_AXI_04_WDATA_PARITY),
    .AXI_04_RDATA_PARITY(instHbm_AXI_04_RDATA_PARITY),
    .AXI_05_ACLK(instHbm_AXI_05_ACLK),
    .AXI_05_ARESET_N(instHbm_AXI_05_ARESET_N),
    .AXI_05_ARADDR(instHbm_AXI_05_ARADDR),
    .AXI_05_ARBURST(instHbm_AXI_05_ARBURST),
    .AXI_05_ARID(instHbm_AXI_05_ARID),
    .AXI_05_ARLEN(instHbm_AXI_05_ARLEN),
    .AXI_05_ARSIZE(instHbm_AXI_05_ARSIZE),
    .AXI_05_ARVALID(instHbm_AXI_05_ARVALID),
    .AXI_05_ARREADY(instHbm_AXI_05_ARREADY),
    .AXI_05_AWADDR(instHbm_AXI_05_AWADDR),
    .AXI_05_AWBURST(instHbm_AXI_05_AWBURST),
    .AXI_05_AWID(instHbm_AXI_05_AWID),
    .AXI_05_AWLEN(instHbm_AXI_05_AWLEN),
    .AXI_05_AWSIZE(instHbm_AXI_05_AWSIZE),
    .AXI_05_AWVALID(instHbm_AXI_05_AWVALID),
    .AXI_05_AWREADY(instHbm_AXI_05_AWREADY),
    .AXI_05_WDATA(instHbm_AXI_05_WDATA),
    .AXI_05_WLAST(instHbm_AXI_05_WLAST),
    .AXI_05_WSTRB(instHbm_AXI_05_WSTRB),
    .AXI_05_WVALID(instHbm_AXI_05_WVALID),
    .AXI_05_WREADY(instHbm_AXI_05_WREADY),
    .AXI_05_RDATA(instHbm_AXI_05_RDATA),
    .AXI_05_RID(instHbm_AXI_05_RID),
    .AXI_05_RLAST(instHbm_AXI_05_RLAST),
    .AXI_05_RRESP(instHbm_AXI_05_RRESP),
    .AXI_05_RVALID(instHbm_AXI_05_RVALID),
    .AXI_05_RREADY(instHbm_AXI_05_RREADY),
    .AXI_05_BID(instHbm_AXI_05_BID),
    .AXI_05_BRESP(instHbm_AXI_05_BRESP),
    .AXI_05_BVALID(instHbm_AXI_05_BVALID),
    .AXI_05_BREADY(instHbm_AXI_05_BREADY),
    .AXI_05_WDATA_PARITY(instHbm_AXI_05_WDATA_PARITY),
    .AXI_05_RDATA_PARITY(instHbm_AXI_05_RDATA_PARITY),
    .AXI_06_ACLK(instHbm_AXI_06_ACLK),
    .AXI_06_ARESET_N(instHbm_AXI_06_ARESET_N),
    .AXI_06_ARADDR(instHbm_AXI_06_ARADDR),
    .AXI_06_ARBURST(instHbm_AXI_06_ARBURST),
    .AXI_06_ARID(instHbm_AXI_06_ARID),
    .AXI_06_ARLEN(instHbm_AXI_06_ARLEN),
    .AXI_06_ARSIZE(instHbm_AXI_06_ARSIZE),
    .AXI_06_ARVALID(instHbm_AXI_06_ARVALID),
    .AXI_06_ARREADY(instHbm_AXI_06_ARREADY),
    .AXI_06_AWADDR(instHbm_AXI_06_AWADDR),
    .AXI_06_AWBURST(instHbm_AXI_06_AWBURST),
    .AXI_06_AWID(instHbm_AXI_06_AWID),
    .AXI_06_AWLEN(instHbm_AXI_06_AWLEN),
    .AXI_06_AWSIZE(instHbm_AXI_06_AWSIZE),
    .AXI_06_AWVALID(instHbm_AXI_06_AWVALID),
    .AXI_06_AWREADY(instHbm_AXI_06_AWREADY),
    .AXI_06_WDATA(instHbm_AXI_06_WDATA),
    .AXI_06_WLAST(instHbm_AXI_06_WLAST),
    .AXI_06_WSTRB(instHbm_AXI_06_WSTRB),
    .AXI_06_WVALID(instHbm_AXI_06_WVALID),
    .AXI_06_WREADY(instHbm_AXI_06_WREADY),
    .AXI_06_RDATA(instHbm_AXI_06_RDATA),
    .AXI_06_RID(instHbm_AXI_06_RID),
    .AXI_06_RLAST(instHbm_AXI_06_RLAST),
    .AXI_06_RRESP(instHbm_AXI_06_RRESP),
    .AXI_06_RVALID(instHbm_AXI_06_RVALID),
    .AXI_06_RREADY(instHbm_AXI_06_RREADY),
    .AXI_06_BID(instHbm_AXI_06_BID),
    .AXI_06_BRESP(instHbm_AXI_06_BRESP),
    .AXI_06_BVALID(instHbm_AXI_06_BVALID),
    .AXI_06_BREADY(instHbm_AXI_06_BREADY),
    .AXI_06_WDATA_PARITY(instHbm_AXI_06_WDATA_PARITY),
    .AXI_06_RDATA_PARITY(instHbm_AXI_06_RDATA_PARITY),
    .AXI_07_ACLK(instHbm_AXI_07_ACLK),
    .AXI_07_ARESET_N(instHbm_AXI_07_ARESET_N),
    .AXI_07_ARADDR(instHbm_AXI_07_ARADDR),
    .AXI_07_ARBURST(instHbm_AXI_07_ARBURST),
    .AXI_07_ARID(instHbm_AXI_07_ARID),
    .AXI_07_ARLEN(instHbm_AXI_07_ARLEN),
    .AXI_07_ARSIZE(instHbm_AXI_07_ARSIZE),
    .AXI_07_ARVALID(instHbm_AXI_07_ARVALID),
    .AXI_07_ARREADY(instHbm_AXI_07_ARREADY),
    .AXI_07_AWADDR(instHbm_AXI_07_AWADDR),
    .AXI_07_AWBURST(instHbm_AXI_07_AWBURST),
    .AXI_07_AWID(instHbm_AXI_07_AWID),
    .AXI_07_AWLEN(instHbm_AXI_07_AWLEN),
    .AXI_07_AWSIZE(instHbm_AXI_07_AWSIZE),
    .AXI_07_AWVALID(instHbm_AXI_07_AWVALID),
    .AXI_07_AWREADY(instHbm_AXI_07_AWREADY),
    .AXI_07_WDATA(instHbm_AXI_07_WDATA),
    .AXI_07_WLAST(instHbm_AXI_07_WLAST),
    .AXI_07_WSTRB(instHbm_AXI_07_WSTRB),
    .AXI_07_WVALID(instHbm_AXI_07_WVALID),
    .AXI_07_WREADY(instHbm_AXI_07_WREADY),
    .AXI_07_RDATA(instHbm_AXI_07_RDATA),
    .AXI_07_RID(instHbm_AXI_07_RID),
    .AXI_07_RLAST(instHbm_AXI_07_RLAST),
    .AXI_07_RRESP(instHbm_AXI_07_RRESP),
    .AXI_07_RVALID(instHbm_AXI_07_RVALID),
    .AXI_07_RREADY(instHbm_AXI_07_RREADY),
    .AXI_07_BID(instHbm_AXI_07_BID),
    .AXI_07_BRESP(instHbm_AXI_07_BRESP),
    .AXI_07_BVALID(instHbm_AXI_07_BVALID),
    .AXI_07_BREADY(instHbm_AXI_07_BREADY),
    .AXI_07_WDATA_PARITY(instHbm_AXI_07_WDATA_PARITY),
    .AXI_07_RDATA_PARITY(instHbm_AXI_07_RDATA_PARITY),
    .AXI_08_ACLK(instHbm_AXI_08_ACLK),
    .AXI_08_ARESET_N(instHbm_AXI_08_ARESET_N),
    .AXI_08_ARADDR(instHbm_AXI_08_ARADDR),
    .AXI_08_ARBURST(instHbm_AXI_08_ARBURST),
    .AXI_08_ARID(instHbm_AXI_08_ARID),
    .AXI_08_ARLEN(instHbm_AXI_08_ARLEN),
    .AXI_08_ARSIZE(instHbm_AXI_08_ARSIZE),
    .AXI_08_ARVALID(instHbm_AXI_08_ARVALID),
    .AXI_08_ARREADY(instHbm_AXI_08_ARREADY),
    .AXI_08_AWADDR(instHbm_AXI_08_AWADDR),
    .AXI_08_AWBURST(instHbm_AXI_08_AWBURST),
    .AXI_08_AWID(instHbm_AXI_08_AWID),
    .AXI_08_AWLEN(instHbm_AXI_08_AWLEN),
    .AXI_08_AWSIZE(instHbm_AXI_08_AWSIZE),
    .AXI_08_AWVALID(instHbm_AXI_08_AWVALID),
    .AXI_08_AWREADY(instHbm_AXI_08_AWREADY),
    .AXI_08_WDATA(instHbm_AXI_08_WDATA),
    .AXI_08_WLAST(instHbm_AXI_08_WLAST),
    .AXI_08_WSTRB(instHbm_AXI_08_WSTRB),
    .AXI_08_WVALID(instHbm_AXI_08_WVALID),
    .AXI_08_WREADY(instHbm_AXI_08_WREADY),
    .AXI_08_RDATA(instHbm_AXI_08_RDATA),
    .AXI_08_RID(instHbm_AXI_08_RID),
    .AXI_08_RLAST(instHbm_AXI_08_RLAST),
    .AXI_08_RRESP(instHbm_AXI_08_RRESP),
    .AXI_08_RVALID(instHbm_AXI_08_RVALID),
    .AXI_08_RREADY(instHbm_AXI_08_RREADY),
    .AXI_08_BID(instHbm_AXI_08_BID),
    .AXI_08_BRESP(instHbm_AXI_08_BRESP),
    .AXI_08_BVALID(instHbm_AXI_08_BVALID),
    .AXI_08_BREADY(instHbm_AXI_08_BREADY),
    .AXI_08_WDATA_PARITY(instHbm_AXI_08_WDATA_PARITY),
    .AXI_08_RDATA_PARITY(instHbm_AXI_08_RDATA_PARITY),
    .AXI_09_ACLK(instHbm_AXI_09_ACLK),
    .AXI_09_ARESET_N(instHbm_AXI_09_ARESET_N),
    .AXI_09_ARADDR(instHbm_AXI_09_ARADDR),
    .AXI_09_ARBURST(instHbm_AXI_09_ARBURST),
    .AXI_09_ARID(instHbm_AXI_09_ARID),
    .AXI_09_ARLEN(instHbm_AXI_09_ARLEN),
    .AXI_09_ARSIZE(instHbm_AXI_09_ARSIZE),
    .AXI_09_ARVALID(instHbm_AXI_09_ARVALID),
    .AXI_09_ARREADY(instHbm_AXI_09_ARREADY),
    .AXI_09_AWADDR(instHbm_AXI_09_AWADDR),
    .AXI_09_AWBURST(instHbm_AXI_09_AWBURST),
    .AXI_09_AWID(instHbm_AXI_09_AWID),
    .AXI_09_AWLEN(instHbm_AXI_09_AWLEN),
    .AXI_09_AWSIZE(instHbm_AXI_09_AWSIZE),
    .AXI_09_AWVALID(instHbm_AXI_09_AWVALID),
    .AXI_09_AWREADY(instHbm_AXI_09_AWREADY),
    .AXI_09_WDATA(instHbm_AXI_09_WDATA),
    .AXI_09_WLAST(instHbm_AXI_09_WLAST),
    .AXI_09_WSTRB(instHbm_AXI_09_WSTRB),
    .AXI_09_WVALID(instHbm_AXI_09_WVALID),
    .AXI_09_WREADY(instHbm_AXI_09_WREADY),
    .AXI_09_RDATA(instHbm_AXI_09_RDATA),
    .AXI_09_RID(instHbm_AXI_09_RID),
    .AXI_09_RLAST(instHbm_AXI_09_RLAST),
    .AXI_09_RRESP(instHbm_AXI_09_RRESP),
    .AXI_09_RVALID(instHbm_AXI_09_RVALID),
    .AXI_09_RREADY(instHbm_AXI_09_RREADY),
    .AXI_09_BID(instHbm_AXI_09_BID),
    .AXI_09_BRESP(instHbm_AXI_09_BRESP),
    .AXI_09_BVALID(instHbm_AXI_09_BVALID),
    .AXI_09_BREADY(instHbm_AXI_09_BREADY),
    .AXI_09_WDATA_PARITY(instHbm_AXI_09_WDATA_PARITY),
    .AXI_09_RDATA_PARITY(instHbm_AXI_09_RDATA_PARITY),
    .AXI_10_ACLK(instHbm_AXI_10_ACLK),
    .AXI_10_ARESET_N(instHbm_AXI_10_ARESET_N),
    .AXI_10_ARADDR(instHbm_AXI_10_ARADDR),
    .AXI_10_ARBURST(instHbm_AXI_10_ARBURST),
    .AXI_10_ARID(instHbm_AXI_10_ARID),
    .AXI_10_ARLEN(instHbm_AXI_10_ARLEN),
    .AXI_10_ARSIZE(instHbm_AXI_10_ARSIZE),
    .AXI_10_ARVALID(instHbm_AXI_10_ARVALID),
    .AXI_10_ARREADY(instHbm_AXI_10_ARREADY),
    .AXI_10_AWADDR(instHbm_AXI_10_AWADDR),
    .AXI_10_AWBURST(instHbm_AXI_10_AWBURST),
    .AXI_10_AWID(instHbm_AXI_10_AWID),
    .AXI_10_AWLEN(instHbm_AXI_10_AWLEN),
    .AXI_10_AWSIZE(instHbm_AXI_10_AWSIZE),
    .AXI_10_AWVALID(instHbm_AXI_10_AWVALID),
    .AXI_10_AWREADY(instHbm_AXI_10_AWREADY),
    .AXI_10_WDATA(instHbm_AXI_10_WDATA),
    .AXI_10_WLAST(instHbm_AXI_10_WLAST),
    .AXI_10_WSTRB(instHbm_AXI_10_WSTRB),
    .AXI_10_WVALID(instHbm_AXI_10_WVALID),
    .AXI_10_WREADY(instHbm_AXI_10_WREADY),
    .AXI_10_RDATA(instHbm_AXI_10_RDATA),
    .AXI_10_RID(instHbm_AXI_10_RID),
    .AXI_10_RLAST(instHbm_AXI_10_RLAST),
    .AXI_10_RRESP(instHbm_AXI_10_RRESP),
    .AXI_10_RVALID(instHbm_AXI_10_RVALID),
    .AXI_10_RREADY(instHbm_AXI_10_RREADY),
    .AXI_10_BID(instHbm_AXI_10_BID),
    .AXI_10_BRESP(instHbm_AXI_10_BRESP),
    .AXI_10_BVALID(instHbm_AXI_10_BVALID),
    .AXI_10_BREADY(instHbm_AXI_10_BREADY),
    .AXI_10_WDATA_PARITY(instHbm_AXI_10_WDATA_PARITY),
    .AXI_10_RDATA_PARITY(instHbm_AXI_10_RDATA_PARITY),
    .AXI_11_ACLK(instHbm_AXI_11_ACLK),
    .AXI_11_ARESET_N(instHbm_AXI_11_ARESET_N),
    .AXI_11_ARADDR(instHbm_AXI_11_ARADDR),
    .AXI_11_ARBURST(instHbm_AXI_11_ARBURST),
    .AXI_11_ARID(instHbm_AXI_11_ARID),
    .AXI_11_ARLEN(instHbm_AXI_11_ARLEN),
    .AXI_11_ARSIZE(instHbm_AXI_11_ARSIZE),
    .AXI_11_ARVALID(instHbm_AXI_11_ARVALID),
    .AXI_11_ARREADY(instHbm_AXI_11_ARREADY),
    .AXI_11_AWADDR(instHbm_AXI_11_AWADDR),
    .AXI_11_AWBURST(instHbm_AXI_11_AWBURST),
    .AXI_11_AWID(instHbm_AXI_11_AWID),
    .AXI_11_AWLEN(instHbm_AXI_11_AWLEN),
    .AXI_11_AWSIZE(instHbm_AXI_11_AWSIZE),
    .AXI_11_AWVALID(instHbm_AXI_11_AWVALID),
    .AXI_11_AWREADY(instHbm_AXI_11_AWREADY),
    .AXI_11_WDATA(instHbm_AXI_11_WDATA),
    .AXI_11_WLAST(instHbm_AXI_11_WLAST),
    .AXI_11_WSTRB(instHbm_AXI_11_WSTRB),
    .AXI_11_WVALID(instHbm_AXI_11_WVALID),
    .AXI_11_WREADY(instHbm_AXI_11_WREADY),
    .AXI_11_RDATA(instHbm_AXI_11_RDATA),
    .AXI_11_RID(instHbm_AXI_11_RID),
    .AXI_11_RLAST(instHbm_AXI_11_RLAST),
    .AXI_11_RRESP(instHbm_AXI_11_RRESP),
    .AXI_11_RVALID(instHbm_AXI_11_RVALID),
    .AXI_11_RREADY(instHbm_AXI_11_RREADY),
    .AXI_11_BID(instHbm_AXI_11_BID),
    .AXI_11_BRESP(instHbm_AXI_11_BRESP),
    .AXI_11_BVALID(instHbm_AXI_11_BVALID),
    .AXI_11_BREADY(instHbm_AXI_11_BREADY),
    .AXI_11_WDATA_PARITY(instHbm_AXI_11_WDATA_PARITY),
    .AXI_11_RDATA_PARITY(instHbm_AXI_11_RDATA_PARITY),
    .AXI_12_ACLK(instHbm_AXI_12_ACLK),
    .AXI_12_ARESET_N(instHbm_AXI_12_ARESET_N),
    .AXI_12_ARADDR(instHbm_AXI_12_ARADDR),
    .AXI_12_ARBURST(instHbm_AXI_12_ARBURST),
    .AXI_12_ARID(instHbm_AXI_12_ARID),
    .AXI_12_ARLEN(instHbm_AXI_12_ARLEN),
    .AXI_12_ARSIZE(instHbm_AXI_12_ARSIZE),
    .AXI_12_ARVALID(instHbm_AXI_12_ARVALID),
    .AXI_12_ARREADY(instHbm_AXI_12_ARREADY),
    .AXI_12_AWADDR(instHbm_AXI_12_AWADDR),
    .AXI_12_AWBURST(instHbm_AXI_12_AWBURST),
    .AXI_12_AWID(instHbm_AXI_12_AWID),
    .AXI_12_AWLEN(instHbm_AXI_12_AWLEN),
    .AXI_12_AWSIZE(instHbm_AXI_12_AWSIZE),
    .AXI_12_AWVALID(instHbm_AXI_12_AWVALID),
    .AXI_12_AWREADY(instHbm_AXI_12_AWREADY),
    .AXI_12_WDATA(instHbm_AXI_12_WDATA),
    .AXI_12_WLAST(instHbm_AXI_12_WLAST),
    .AXI_12_WSTRB(instHbm_AXI_12_WSTRB),
    .AXI_12_WVALID(instHbm_AXI_12_WVALID),
    .AXI_12_WREADY(instHbm_AXI_12_WREADY),
    .AXI_12_RDATA(instHbm_AXI_12_RDATA),
    .AXI_12_RID(instHbm_AXI_12_RID),
    .AXI_12_RLAST(instHbm_AXI_12_RLAST),
    .AXI_12_RRESP(instHbm_AXI_12_RRESP),
    .AXI_12_RVALID(instHbm_AXI_12_RVALID),
    .AXI_12_RREADY(instHbm_AXI_12_RREADY),
    .AXI_12_BID(instHbm_AXI_12_BID),
    .AXI_12_BRESP(instHbm_AXI_12_BRESP),
    .AXI_12_BVALID(instHbm_AXI_12_BVALID),
    .AXI_12_BREADY(instHbm_AXI_12_BREADY),
    .AXI_12_WDATA_PARITY(instHbm_AXI_12_WDATA_PARITY),
    .AXI_12_RDATA_PARITY(instHbm_AXI_12_RDATA_PARITY),
    .AXI_13_ACLK(instHbm_AXI_13_ACLK),
    .AXI_13_ARESET_N(instHbm_AXI_13_ARESET_N),
    .AXI_13_ARADDR(instHbm_AXI_13_ARADDR),
    .AXI_13_ARBURST(instHbm_AXI_13_ARBURST),
    .AXI_13_ARID(instHbm_AXI_13_ARID),
    .AXI_13_ARLEN(instHbm_AXI_13_ARLEN),
    .AXI_13_ARSIZE(instHbm_AXI_13_ARSIZE),
    .AXI_13_ARVALID(instHbm_AXI_13_ARVALID),
    .AXI_13_ARREADY(instHbm_AXI_13_ARREADY),
    .AXI_13_AWADDR(instHbm_AXI_13_AWADDR),
    .AXI_13_AWBURST(instHbm_AXI_13_AWBURST),
    .AXI_13_AWID(instHbm_AXI_13_AWID),
    .AXI_13_AWLEN(instHbm_AXI_13_AWLEN),
    .AXI_13_AWSIZE(instHbm_AXI_13_AWSIZE),
    .AXI_13_AWVALID(instHbm_AXI_13_AWVALID),
    .AXI_13_AWREADY(instHbm_AXI_13_AWREADY),
    .AXI_13_WDATA(instHbm_AXI_13_WDATA),
    .AXI_13_WLAST(instHbm_AXI_13_WLAST),
    .AXI_13_WSTRB(instHbm_AXI_13_WSTRB),
    .AXI_13_WVALID(instHbm_AXI_13_WVALID),
    .AXI_13_WREADY(instHbm_AXI_13_WREADY),
    .AXI_13_RDATA(instHbm_AXI_13_RDATA),
    .AXI_13_RID(instHbm_AXI_13_RID),
    .AXI_13_RLAST(instHbm_AXI_13_RLAST),
    .AXI_13_RRESP(instHbm_AXI_13_RRESP),
    .AXI_13_RVALID(instHbm_AXI_13_RVALID),
    .AXI_13_RREADY(instHbm_AXI_13_RREADY),
    .AXI_13_BID(instHbm_AXI_13_BID),
    .AXI_13_BRESP(instHbm_AXI_13_BRESP),
    .AXI_13_BVALID(instHbm_AXI_13_BVALID),
    .AXI_13_BREADY(instHbm_AXI_13_BREADY),
    .AXI_13_WDATA_PARITY(instHbm_AXI_13_WDATA_PARITY),
    .AXI_13_RDATA_PARITY(instHbm_AXI_13_RDATA_PARITY),
    .AXI_14_ACLK(instHbm_AXI_14_ACLK),
    .AXI_14_ARESET_N(instHbm_AXI_14_ARESET_N),
    .AXI_14_ARADDR(instHbm_AXI_14_ARADDR),
    .AXI_14_ARBURST(instHbm_AXI_14_ARBURST),
    .AXI_14_ARID(instHbm_AXI_14_ARID),
    .AXI_14_ARLEN(instHbm_AXI_14_ARLEN),
    .AXI_14_ARSIZE(instHbm_AXI_14_ARSIZE),
    .AXI_14_ARVALID(instHbm_AXI_14_ARVALID),
    .AXI_14_ARREADY(instHbm_AXI_14_ARREADY),
    .AXI_14_AWADDR(instHbm_AXI_14_AWADDR),
    .AXI_14_AWBURST(instHbm_AXI_14_AWBURST),
    .AXI_14_AWID(instHbm_AXI_14_AWID),
    .AXI_14_AWLEN(instHbm_AXI_14_AWLEN),
    .AXI_14_AWSIZE(instHbm_AXI_14_AWSIZE),
    .AXI_14_AWVALID(instHbm_AXI_14_AWVALID),
    .AXI_14_AWREADY(instHbm_AXI_14_AWREADY),
    .AXI_14_WDATA(instHbm_AXI_14_WDATA),
    .AXI_14_WLAST(instHbm_AXI_14_WLAST),
    .AXI_14_WSTRB(instHbm_AXI_14_WSTRB),
    .AXI_14_WVALID(instHbm_AXI_14_WVALID),
    .AXI_14_WREADY(instHbm_AXI_14_WREADY),
    .AXI_14_RDATA(instHbm_AXI_14_RDATA),
    .AXI_14_RID(instHbm_AXI_14_RID),
    .AXI_14_RLAST(instHbm_AXI_14_RLAST),
    .AXI_14_RRESP(instHbm_AXI_14_RRESP),
    .AXI_14_RVALID(instHbm_AXI_14_RVALID),
    .AXI_14_RREADY(instHbm_AXI_14_RREADY),
    .AXI_14_BID(instHbm_AXI_14_BID),
    .AXI_14_BRESP(instHbm_AXI_14_BRESP),
    .AXI_14_BVALID(instHbm_AXI_14_BVALID),
    .AXI_14_BREADY(instHbm_AXI_14_BREADY),
    .AXI_14_WDATA_PARITY(instHbm_AXI_14_WDATA_PARITY),
    .AXI_14_RDATA_PARITY(instHbm_AXI_14_RDATA_PARITY),
    .AXI_15_ACLK(instHbm_AXI_15_ACLK),
    .AXI_15_ARESET_N(instHbm_AXI_15_ARESET_N),
    .AXI_15_ARADDR(instHbm_AXI_15_ARADDR),
    .AXI_15_ARBURST(instHbm_AXI_15_ARBURST),
    .AXI_15_ARID(instHbm_AXI_15_ARID),
    .AXI_15_ARLEN(instHbm_AXI_15_ARLEN),
    .AXI_15_ARSIZE(instHbm_AXI_15_ARSIZE),
    .AXI_15_ARVALID(instHbm_AXI_15_ARVALID),
    .AXI_15_ARREADY(instHbm_AXI_15_ARREADY),
    .AXI_15_AWADDR(instHbm_AXI_15_AWADDR),
    .AXI_15_AWBURST(instHbm_AXI_15_AWBURST),
    .AXI_15_AWID(instHbm_AXI_15_AWID),
    .AXI_15_AWLEN(instHbm_AXI_15_AWLEN),
    .AXI_15_AWSIZE(instHbm_AXI_15_AWSIZE),
    .AXI_15_AWVALID(instHbm_AXI_15_AWVALID),
    .AXI_15_AWREADY(instHbm_AXI_15_AWREADY),
    .AXI_15_WDATA(instHbm_AXI_15_WDATA),
    .AXI_15_WLAST(instHbm_AXI_15_WLAST),
    .AXI_15_WSTRB(instHbm_AXI_15_WSTRB),
    .AXI_15_WVALID(instHbm_AXI_15_WVALID),
    .AXI_15_WREADY(instHbm_AXI_15_WREADY),
    .AXI_15_RDATA(instHbm_AXI_15_RDATA),
    .AXI_15_RID(instHbm_AXI_15_RID),
    .AXI_15_RLAST(instHbm_AXI_15_RLAST),
    .AXI_15_RRESP(instHbm_AXI_15_RRESP),
    .AXI_15_RVALID(instHbm_AXI_15_RVALID),
    .AXI_15_RREADY(instHbm_AXI_15_RREADY),
    .AXI_15_BID(instHbm_AXI_15_BID),
    .AXI_15_BRESP(instHbm_AXI_15_BRESP),
    .AXI_15_BVALID(instHbm_AXI_15_BVALID),
    .AXI_15_BREADY(instHbm_AXI_15_BREADY),
    .AXI_15_WDATA_PARITY(instHbm_AXI_15_WDATA_PARITY),
    .AXI_15_RDATA_PARITY(instHbm_AXI_15_RDATA_PARITY),
    .AXI_16_ACLK(instHbm_AXI_16_ACLK),
    .AXI_16_ARESET_N(instHbm_AXI_16_ARESET_N),
    .AXI_16_ARADDR(instHbm_AXI_16_ARADDR),
    .AXI_16_ARBURST(instHbm_AXI_16_ARBURST),
    .AXI_16_ARID(instHbm_AXI_16_ARID),
    .AXI_16_ARLEN(instHbm_AXI_16_ARLEN),
    .AXI_16_ARSIZE(instHbm_AXI_16_ARSIZE),
    .AXI_16_ARVALID(instHbm_AXI_16_ARVALID),
    .AXI_16_ARREADY(instHbm_AXI_16_ARREADY),
    .AXI_16_AWADDR(instHbm_AXI_16_AWADDR),
    .AXI_16_AWBURST(instHbm_AXI_16_AWBURST),
    .AXI_16_AWID(instHbm_AXI_16_AWID),
    .AXI_16_AWLEN(instHbm_AXI_16_AWLEN),
    .AXI_16_AWSIZE(instHbm_AXI_16_AWSIZE),
    .AXI_16_AWVALID(instHbm_AXI_16_AWVALID),
    .AXI_16_AWREADY(instHbm_AXI_16_AWREADY),
    .AXI_16_WDATA(instHbm_AXI_16_WDATA),
    .AXI_16_WLAST(instHbm_AXI_16_WLAST),
    .AXI_16_WSTRB(instHbm_AXI_16_WSTRB),
    .AXI_16_WVALID(instHbm_AXI_16_WVALID),
    .AXI_16_WREADY(instHbm_AXI_16_WREADY),
    .AXI_16_RDATA(instHbm_AXI_16_RDATA),
    .AXI_16_RID(instHbm_AXI_16_RID),
    .AXI_16_RLAST(instHbm_AXI_16_RLAST),
    .AXI_16_RRESP(instHbm_AXI_16_RRESP),
    .AXI_16_RVALID(instHbm_AXI_16_RVALID),
    .AXI_16_RREADY(instHbm_AXI_16_RREADY),
    .AXI_16_BID(instHbm_AXI_16_BID),
    .AXI_16_BRESP(instHbm_AXI_16_BRESP),
    .AXI_16_BVALID(instHbm_AXI_16_BVALID),
    .AXI_16_BREADY(instHbm_AXI_16_BREADY),
    .AXI_16_WDATA_PARITY(instHbm_AXI_16_WDATA_PARITY),
    .AXI_16_RDATA_PARITY(instHbm_AXI_16_RDATA_PARITY),
    .AXI_17_ACLK(instHbm_AXI_17_ACLK),
    .AXI_17_ARESET_N(instHbm_AXI_17_ARESET_N),
    .AXI_17_ARADDR(instHbm_AXI_17_ARADDR),
    .AXI_17_ARBURST(instHbm_AXI_17_ARBURST),
    .AXI_17_ARID(instHbm_AXI_17_ARID),
    .AXI_17_ARLEN(instHbm_AXI_17_ARLEN),
    .AXI_17_ARSIZE(instHbm_AXI_17_ARSIZE),
    .AXI_17_ARVALID(instHbm_AXI_17_ARVALID),
    .AXI_17_ARREADY(instHbm_AXI_17_ARREADY),
    .AXI_17_AWADDR(instHbm_AXI_17_AWADDR),
    .AXI_17_AWBURST(instHbm_AXI_17_AWBURST),
    .AXI_17_AWID(instHbm_AXI_17_AWID),
    .AXI_17_AWLEN(instHbm_AXI_17_AWLEN),
    .AXI_17_AWSIZE(instHbm_AXI_17_AWSIZE),
    .AXI_17_AWVALID(instHbm_AXI_17_AWVALID),
    .AXI_17_AWREADY(instHbm_AXI_17_AWREADY),
    .AXI_17_WDATA(instHbm_AXI_17_WDATA),
    .AXI_17_WLAST(instHbm_AXI_17_WLAST),
    .AXI_17_WSTRB(instHbm_AXI_17_WSTRB),
    .AXI_17_WVALID(instHbm_AXI_17_WVALID),
    .AXI_17_WREADY(instHbm_AXI_17_WREADY),
    .AXI_17_RDATA(instHbm_AXI_17_RDATA),
    .AXI_17_RID(instHbm_AXI_17_RID),
    .AXI_17_RLAST(instHbm_AXI_17_RLAST),
    .AXI_17_RRESP(instHbm_AXI_17_RRESP),
    .AXI_17_RVALID(instHbm_AXI_17_RVALID),
    .AXI_17_RREADY(instHbm_AXI_17_RREADY),
    .AXI_17_BID(instHbm_AXI_17_BID),
    .AXI_17_BRESP(instHbm_AXI_17_BRESP),
    .AXI_17_BVALID(instHbm_AXI_17_BVALID),
    .AXI_17_BREADY(instHbm_AXI_17_BREADY),
    .AXI_17_WDATA_PARITY(instHbm_AXI_17_WDATA_PARITY),
    .AXI_17_RDATA_PARITY(instHbm_AXI_17_RDATA_PARITY),
    .AXI_18_ACLK(instHbm_AXI_18_ACLK),
    .AXI_18_ARESET_N(instHbm_AXI_18_ARESET_N),
    .AXI_18_ARADDR(instHbm_AXI_18_ARADDR),
    .AXI_18_ARBURST(instHbm_AXI_18_ARBURST),
    .AXI_18_ARID(instHbm_AXI_18_ARID),
    .AXI_18_ARLEN(instHbm_AXI_18_ARLEN),
    .AXI_18_ARSIZE(instHbm_AXI_18_ARSIZE),
    .AXI_18_ARVALID(instHbm_AXI_18_ARVALID),
    .AXI_18_ARREADY(instHbm_AXI_18_ARREADY),
    .AXI_18_AWADDR(instHbm_AXI_18_AWADDR),
    .AXI_18_AWBURST(instHbm_AXI_18_AWBURST),
    .AXI_18_AWID(instHbm_AXI_18_AWID),
    .AXI_18_AWLEN(instHbm_AXI_18_AWLEN),
    .AXI_18_AWSIZE(instHbm_AXI_18_AWSIZE),
    .AXI_18_AWVALID(instHbm_AXI_18_AWVALID),
    .AXI_18_AWREADY(instHbm_AXI_18_AWREADY),
    .AXI_18_WDATA(instHbm_AXI_18_WDATA),
    .AXI_18_WLAST(instHbm_AXI_18_WLAST),
    .AXI_18_WSTRB(instHbm_AXI_18_WSTRB),
    .AXI_18_WVALID(instHbm_AXI_18_WVALID),
    .AXI_18_WREADY(instHbm_AXI_18_WREADY),
    .AXI_18_RDATA(instHbm_AXI_18_RDATA),
    .AXI_18_RID(instHbm_AXI_18_RID),
    .AXI_18_RLAST(instHbm_AXI_18_RLAST),
    .AXI_18_RRESP(instHbm_AXI_18_RRESP),
    .AXI_18_RVALID(instHbm_AXI_18_RVALID),
    .AXI_18_RREADY(instHbm_AXI_18_RREADY),
    .AXI_18_BID(instHbm_AXI_18_BID),
    .AXI_18_BRESP(instHbm_AXI_18_BRESP),
    .AXI_18_BVALID(instHbm_AXI_18_BVALID),
    .AXI_18_BREADY(instHbm_AXI_18_BREADY),
    .AXI_18_WDATA_PARITY(instHbm_AXI_18_WDATA_PARITY),
    .AXI_18_RDATA_PARITY(instHbm_AXI_18_RDATA_PARITY),
    .AXI_19_ACLK(instHbm_AXI_19_ACLK),
    .AXI_19_ARESET_N(instHbm_AXI_19_ARESET_N),
    .AXI_19_ARADDR(instHbm_AXI_19_ARADDR),
    .AXI_19_ARBURST(instHbm_AXI_19_ARBURST),
    .AXI_19_ARID(instHbm_AXI_19_ARID),
    .AXI_19_ARLEN(instHbm_AXI_19_ARLEN),
    .AXI_19_ARSIZE(instHbm_AXI_19_ARSIZE),
    .AXI_19_ARVALID(instHbm_AXI_19_ARVALID),
    .AXI_19_ARREADY(instHbm_AXI_19_ARREADY),
    .AXI_19_AWADDR(instHbm_AXI_19_AWADDR),
    .AXI_19_AWBURST(instHbm_AXI_19_AWBURST),
    .AXI_19_AWID(instHbm_AXI_19_AWID),
    .AXI_19_AWLEN(instHbm_AXI_19_AWLEN),
    .AXI_19_AWSIZE(instHbm_AXI_19_AWSIZE),
    .AXI_19_AWVALID(instHbm_AXI_19_AWVALID),
    .AXI_19_AWREADY(instHbm_AXI_19_AWREADY),
    .AXI_19_WDATA(instHbm_AXI_19_WDATA),
    .AXI_19_WLAST(instHbm_AXI_19_WLAST),
    .AXI_19_WSTRB(instHbm_AXI_19_WSTRB),
    .AXI_19_WVALID(instHbm_AXI_19_WVALID),
    .AXI_19_WREADY(instHbm_AXI_19_WREADY),
    .AXI_19_RDATA(instHbm_AXI_19_RDATA),
    .AXI_19_RID(instHbm_AXI_19_RID),
    .AXI_19_RLAST(instHbm_AXI_19_RLAST),
    .AXI_19_RRESP(instHbm_AXI_19_RRESP),
    .AXI_19_RVALID(instHbm_AXI_19_RVALID),
    .AXI_19_RREADY(instHbm_AXI_19_RREADY),
    .AXI_19_BID(instHbm_AXI_19_BID),
    .AXI_19_BRESP(instHbm_AXI_19_BRESP),
    .AXI_19_BVALID(instHbm_AXI_19_BVALID),
    .AXI_19_BREADY(instHbm_AXI_19_BREADY),
    .AXI_19_WDATA_PARITY(instHbm_AXI_19_WDATA_PARITY),
    .AXI_19_RDATA_PARITY(instHbm_AXI_19_RDATA_PARITY),
    .AXI_20_ACLK(instHbm_AXI_20_ACLK),
    .AXI_20_ARESET_N(instHbm_AXI_20_ARESET_N),
    .AXI_20_ARADDR(instHbm_AXI_20_ARADDR),
    .AXI_20_ARBURST(instHbm_AXI_20_ARBURST),
    .AXI_20_ARID(instHbm_AXI_20_ARID),
    .AXI_20_ARLEN(instHbm_AXI_20_ARLEN),
    .AXI_20_ARSIZE(instHbm_AXI_20_ARSIZE),
    .AXI_20_ARVALID(instHbm_AXI_20_ARVALID),
    .AXI_20_ARREADY(instHbm_AXI_20_ARREADY),
    .AXI_20_AWADDR(instHbm_AXI_20_AWADDR),
    .AXI_20_AWBURST(instHbm_AXI_20_AWBURST),
    .AXI_20_AWID(instHbm_AXI_20_AWID),
    .AXI_20_AWLEN(instHbm_AXI_20_AWLEN),
    .AXI_20_AWSIZE(instHbm_AXI_20_AWSIZE),
    .AXI_20_AWVALID(instHbm_AXI_20_AWVALID),
    .AXI_20_AWREADY(instHbm_AXI_20_AWREADY),
    .AXI_20_WDATA(instHbm_AXI_20_WDATA),
    .AXI_20_WLAST(instHbm_AXI_20_WLAST),
    .AXI_20_WSTRB(instHbm_AXI_20_WSTRB),
    .AXI_20_WVALID(instHbm_AXI_20_WVALID),
    .AXI_20_WREADY(instHbm_AXI_20_WREADY),
    .AXI_20_RDATA(instHbm_AXI_20_RDATA),
    .AXI_20_RID(instHbm_AXI_20_RID),
    .AXI_20_RLAST(instHbm_AXI_20_RLAST),
    .AXI_20_RRESP(instHbm_AXI_20_RRESP),
    .AXI_20_RVALID(instHbm_AXI_20_RVALID),
    .AXI_20_RREADY(instHbm_AXI_20_RREADY),
    .AXI_20_BID(instHbm_AXI_20_BID),
    .AXI_20_BRESP(instHbm_AXI_20_BRESP),
    .AXI_20_BVALID(instHbm_AXI_20_BVALID),
    .AXI_20_BREADY(instHbm_AXI_20_BREADY),
    .AXI_20_WDATA_PARITY(instHbm_AXI_20_WDATA_PARITY),
    .AXI_20_RDATA_PARITY(instHbm_AXI_20_RDATA_PARITY),
    .AXI_21_ACLK(instHbm_AXI_21_ACLK),
    .AXI_21_ARESET_N(instHbm_AXI_21_ARESET_N),
    .AXI_21_ARADDR(instHbm_AXI_21_ARADDR),
    .AXI_21_ARBURST(instHbm_AXI_21_ARBURST),
    .AXI_21_ARID(instHbm_AXI_21_ARID),
    .AXI_21_ARLEN(instHbm_AXI_21_ARLEN),
    .AXI_21_ARSIZE(instHbm_AXI_21_ARSIZE),
    .AXI_21_ARVALID(instHbm_AXI_21_ARVALID),
    .AXI_21_ARREADY(instHbm_AXI_21_ARREADY),
    .AXI_21_AWADDR(instHbm_AXI_21_AWADDR),
    .AXI_21_AWBURST(instHbm_AXI_21_AWBURST),
    .AXI_21_AWID(instHbm_AXI_21_AWID),
    .AXI_21_AWLEN(instHbm_AXI_21_AWLEN),
    .AXI_21_AWSIZE(instHbm_AXI_21_AWSIZE),
    .AXI_21_AWVALID(instHbm_AXI_21_AWVALID),
    .AXI_21_AWREADY(instHbm_AXI_21_AWREADY),
    .AXI_21_WDATA(instHbm_AXI_21_WDATA),
    .AXI_21_WLAST(instHbm_AXI_21_WLAST),
    .AXI_21_WSTRB(instHbm_AXI_21_WSTRB),
    .AXI_21_WVALID(instHbm_AXI_21_WVALID),
    .AXI_21_WREADY(instHbm_AXI_21_WREADY),
    .AXI_21_RDATA(instHbm_AXI_21_RDATA),
    .AXI_21_RID(instHbm_AXI_21_RID),
    .AXI_21_RLAST(instHbm_AXI_21_RLAST),
    .AXI_21_RRESP(instHbm_AXI_21_RRESP),
    .AXI_21_RVALID(instHbm_AXI_21_RVALID),
    .AXI_21_RREADY(instHbm_AXI_21_RREADY),
    .AXI_21_BID(instHbm_AXI_21_BID),
    .AXI_21_BRESP(instHbm_AXI_21_BRESP),
    .AXI_21_BVALID(instHbm_AXI_21_BVALID),
    .AXI_21_BREADY(instHbm_AXI_21_BREADY),
    .AXI_21_WDATA_PARITY(instHbm_AXI_21_WDATA_PARITY),
    .AXI_21_RDATA_PARITY(instHbm_AXI_21_RDATA_PARITY),
    .AXI_22_ACLK(instHbm_AXI_22_ACLK),
    .AXI_22_ARESET_N(instHbm_AXI_22_ARESET_N),
    .AXI_22_ARADDR(instHbm_AXI_22_ARADDR),
    .AXI_22_ARBURST(instHbm_AXI_22_ARBURST),
    .AXI_22_ARID(instHbm_AXI_22_ARID),
    .AXI_22_ARLEN(instHbm_AXI_22_ARLEN),
    .AXI_22_ARSIZE(instHbm_AXI_22_ARSIZE),
    .AXI_22_ARVALID(instHbm_AXI_22_ARVALID),
    .AXI_22_ARREADY(instHbm_AXI_22_ARREADY),
    .AXI_22_AWADDR(instHbm_AXI_22_AWADDR),
    .AXI_22_AWBURST(instHbm_AXI_22_AWBURST),
    .AXI_22_AWID(instHbm_AXI_22_AWID),
    .AXI_22_AWLEN(instHbm_AXI_22_AWLEN),
    .AXI_22_AWSIZE(instHbm_AXI_22_AWSIZE),
    .AXI_22_AWVALID(instHbm_AXI_22_AWVALID),
    .AXI_22_AWREADY(instHbm_AXI_22_AWREADY),
    .AXI_22_WDATA(instHbm_AXI_22_WDATA),
    .AXI_22_WLAST(instHbm_AXI_22_WLAST),
    .AXI_22_WSTRB(instHbm_AXI_22_WSTRB),
    .AXI_22_WVALID(instHbm_AXI_22_WVALID),
    .AXI_22_WREADY(instHbm_AXI_22_WREADY),
    .AXI_22_RDATA(instHbm_AXI_22_RDATA),
    .AXI_22_RID(instHbm_AXI_22_RID),
    .AXI_22_RLAST(instHbm_AXI_22_RLAST),
    .AXI_22_RRESP(instHbm_AXI_22_RRESP),
    .AXI_22_RVALID(instHbm_AXI_22_RVALID),
    .AXI_22_RREADY(instHbm_AXI_22_RREADY),
    .AXI_22_BID(instHbm_AXI_22_BID),
    .AXI_22_BRESP(instHbm_AXI_22_BRESP),
    .AXI_22_BVALID(instHbm_AXI_22_BVALID),
    .AXI_22_BREADY(instHbm_AXI_22_BREADY),
    .AXI_22_WDATA_PARITY(instHbm_AXI_22_WDATA_PARITY),
    .AXI_22_RDATA_PARITY(instHbm_AXI_22_RDATA_PARITY),
    .AXI_23_ACLK(instHbm_AXI_23_ACLK),
    .AXI_23_ARESET_N(instHbm_AXI_23_ARESET_N),
    .AXI_23_ARADDR(instHbm_AXI_23_ARADDR),
    .AXI_23_ARBURST(instHbm_AXI_23_ARBURST),
    .AXI_23_ARID(instHbm_AXI_23_ARID),
    .AXI_23_ARLEN(instHbm_AXI_23_ARLEN),
    .AXI_23_ARSIZE(instHbm_AXI_23_ARSIZE),
    .AXI_23_ARVALID(instHbm_AXI_23_ARVALID),
    .AXI_23_ARREADY(instHbm_AXI_23_ARREADY),
    .AXI_23_AWADDR(instHbm_AXI_23_AWADDR),
    .AXI_23_AWBURST(instHbm_AXI_23_AWBURST),
    .AXI_23_AWID(instHbm_AXI_23_AWID),
    .AXI_23_AWLEN(instHbm_AXI_23_AWLEN),
    .AXI_23_AWSIZE(instHbm_AXI_23_AWSIZE),
    .AXI_23_AWVALID(instHbm_AXI_23_AWVALID),
    .AXI_23_AWREADY(instHbm_AXI_23_AWREADY),
    .AXI_23_WDATA(instHbm_AXI_23_WDATA),
    .AXI_23_WLAST(instHbm_AXI_23_WLAST),
    .AXI_23_WSTRB(instHbm_AXI_23_WSTRB),
    .AXI_23_WVALID(instHbm_AXI_23_WVALID),
    .AXI_23_WREADY(instHbm_AXI_23_WREADY),
    .AXI_23_RDATA(instHbm_AXI_23_RDATA),
    .AXI_23_RID(instHbm_AXI_23_RID),
    .AXI_23_RLAST(instHbm_AXI_23_RLAST),
    .AXI_23_RRESP(instHbm_AXI_23_RRESP),
    .AXI_23_RVALID(instHbm_AXI_23_RVALID),
    .AXI_23_RREADY(instHbm_AXI_23_RREADY),
    .AXI_23_BID(instHbm_AXI_23_BID),
    .AXI_23_BRESP(instHbm_AXI_23_BRESP),
    .AXI_23_BVALID(instHbm_AXI_23_BVALID),
    .AXI_23_BREADY(instHbm_AXI_23_BREADY),
    .AXI_23_WDATA_PARITY(instHbm_AXI_23_WDATA_PARITY),
    .AXI_23_RDATA_PARITY(instHbm_AXI_23_RDATA_PARITY),
    .AXI_24_ACLK(instHbm_AXI_24_ACLK),
    .AXI_24_ARESET_N(instHbm_AXI_24_ARESET_N),
    .AXI_24_ARADDR(instHbm_AXI_24_ARADDR),
    .AXI_24_ARBURST(instHbm_AXI_24_ARBURST),
    .AXI_24_ARID(instHbm_AXI_24_ARID),
    .AXI_24_ARLEN(instHbm_AXI_24_ARLEN),
    .AXI_24_ARSIZE(instHbm_AXI_24_ARSIZE),
    .AXI_24_ARVALID(instHbm_AXI_24_ARVALID),
    .AXI_24_ARREADY(instHbm_AXI_24_ARREADY),
    .AXI_24_AWADDR(instHbm_AXI_24_AWADDR),
    .AXI_24_AWBURST(instHbm_AXI_24_AWBURST),
    .AXI_24_AWID(instHbm_AXI_24_AWID),
    .AXI_24_AWLEN(instHbm_AXI_24_AWLEN),
    .AXI_24_AWSIZE(instHbm_AXI_24_AWSIZE),
    .AXI_24_AWVALID(instHbm_AXI_24_AWVALID),
    .AXI_24_AWREADY(instHbm_AXI_24_AWREADY),
    .AXI_24_WDATA(instHbm_AXI_24_WDATA),
    .AXI_24_WLAST(instHbm_AXI_24_WLAST),
    .AXI_24_WSTRB(instHbm_AXI_24_WSTRB),
    .AXI_24_WVALID(instHbm_AXI_24_WVALID),
    .AXI_24_WREADY(instHbm_AXI_24_WREADY),
    .AXI_24_RDATA(instHbm_AXI_24_RDATA),
    .AXI_24_RID(instHbm_AXI_24_RID),
    .AXI_24_RLAST(instHbm_AXI_24_RLAST),
    .AXI_24_RRESP(instHbm_AXI_24_RRESP),
    .AXI_24_RVALID(instHbm_AXI_24_RVALID),
    .AXI_24_RREADY(instHbm_AXI_24_RREADY),
    .AXI_24_BID(instHbm_AXI_24_BID),
    .AXI_24_BRESP(instHbm_AXI_24_BRESP),
    .AXI_24_BVALID(instHbm_AXI_24_BVALID),
    .AXI_24_BREADY(instHbm_AXI_24_BREADY),
    .AXI_24_WDATA_PARITY(instHbm_AXI_24_WDATA_PARITY),
    .AXI_24_RDATA_PARITY(instHbm_AXI_24_RDATA_PARITY),
    .AXI_25_ACLK(instHbm_AXI_25_ACLK),
    .AXI_25_ARESET_N(instHbm_AXI_25_ARESET_N),
    .AXI_25_ARADDR(instHbm_AXI_25_ARADDR),
    .AXI_25_ARBURST(instHbm_AXI_25_ARBURST),
    .AXI_25_ARID(instHbm_AXI_25_ARID),
    .AXI_25_ARLEN(instHbm_AXI_25_ARLEN),
    .AXI_25_ARSIZE(instHbm_AXI_25_ARSIZE),
    .AXI_25_ARVALID(instHbm_AXI_25_ARVALID),
    .AXI_25_ARREADY(instHbm_AXI_25_ARREADY),
    .AXI_25_AWADDR(instHbm_AXI_25_AWADDR),
    .AXI_25_AWBURST(instHbm_AXI_25_AWBURST),
    .AXI_25_AWID(instHbm_AXI_25_AWID),
    .AXI_25_AWLEN(instHbm_AXI_25_AWLEN),
    .AXI_25_AWSIZE(instHbm_AXI_25_AWSIZE),
    .AXI_25_AWVALID(instHbm_AXI_25_AWVALID),
    .AXI_25_AWREADY(instHbm_AXI_25_AWREADY),
    .AXI_25_WDATA(instHbm_AXI_25_WDATA),
    .AXI_25_WLAST(instHbm_AXI_25_WLAST),
    .AXI_25_WSTRB(instHbm_AXI_25_WSTRB),
    .AXI_25_WVALID(instHbm_AXI_25_WVALID),
    .AXI_25_WREADY(instHbm_AXI_25_WREADY),
    .AXI_25_RDATA(instHbm_AXI_25_RDATA),
    .AXI_25_RID(instHbm_AXI_25_RID),
    .AXI_25_RLAST(instHbm_AXI_25_RLAST),
    .AXI_25_RRESP(instHbm_AXI_25_RRESP),
    .AXI_25_RVALID(instHbm_AXI_25_RVALID),
    .AXI_25_RREADY(instHbm_AXI_25_RREADY),
    .AXI_25_BID(instHbm_AXI_25_BID),
    .AXI_25_BRESP(instHbm_AXI_25_BRESP),
    .AXI_25_BVALID(instHbm_AXI_25_BVALID),
    .AXI_25_BREADY(instHbm_AXI_25_BREADY),
    .AXI_25_WDATA_PARITY(instHbm_AXI_25_WDATA_PARITY),
    .AXI_25_RDATA_PARITY(instHbm_AXI_25_RDATA_PARITY),
    .AXI_26_ACLK(instHbm_AXI_26_ACLK),
    .AXI_26_ARESET_N(instHbm_AXI_26_ARESET_N),
    .AXI_26_ARADDR(instHbm_AXI_26_ARADDR),
    .AXI_26_ARBURST(instHbm_AXI_26_ARBURST),
    .AXI_26_ARID(instHbm_AXI_26_ARID),
    .AXI_26_ARLEN(instHbm_AXI_26_ARLEN),
    .AXI_26_ARSIZE(instHbm_AXI_26_ARSIZE),
    .AXI_26_ARVALID(instHbm_AXI_26_ARVALID),
    .AXI_26_ARREADY(instHbm_AXI_26_ARREADY),
    .AXI_26_AWADDR(instHbm_AXI_26_AWADDR),
    .AXI_26_AWBURST(instHbm_AXI_26_AWBURST),
    .AXI_26_AWID(instHbm_AXI_26_AWID),
    .AXI_26_AWLEN(instHbm_AXI_26_AWLEN),
    .AXI_26_AWSIZE(instHbm_AXI_26_AWSIZE),
    .AXI_26_AWVALID(instHbm_AXI_26_AWVALID),
    .AXI_26_AWREADY(instHbm_AXI_26_AWREADY),
    .AXI_26_WDATA(instHbm_AXI_26_WDATA),
    .AXI_26_WLAST(instHbm_AXI_26_WLAST),
    .AXI_26_WSTRB(instHbm_AXI_26_WSTRB),
    .AXI_26_WVALID(instHbm_AXI_26_WVALID),
    .AXI_26_WREADY(instHbm_AXI_26_WREADY),
    .AXI_26_RDATA(instHbm_AXI_26_RDATA),
    .AXI_26_RID(instHbm_AXI_26_RID),
    .AXI_26_RLAST(instHbm_AXI_26_RLAST),
    .AXI_26_RRESP(instHbm_AXI_26_RRESP),
    .AXI_26_RVALID(instHbm_AXI_26_RVALID),
    .AXI_26_RREADY(instHbm_AXI_26_RREADY),
    .AXI_26_BID(instHbm_AXI_26_BID),
    .AXI_26_BRESP(instHbm_AXI_26_BRESP),
    .AXI_26_BVALID(instHbm_AXI_26_BVALID),
    .AXI_26_BREADY(instHbm_AXI_26_BREADY),
    .AXI_26_WDATA_PARITY(instHbm_AXI_26_WDATA_PARITY),
    .AXI_26_RDATA_PARITY(instHbm_AXI_26_RDATA_PARITY),
    .AXI_27_ACLK(instHbm_AXI_27_ACLK),
    .AXI_27_ARESET_N(instHbm_AXI_27_ARESET_N),
    .AXI_27_ARADDR(instHbm_AXI_27_ARADDR),
    .AXI_27_ARBURST(instHbm_AXI_27_ARBURST),
    .AXI_27_ARID(instHbm_AXI_27_ARID),
    .AXI_27_ARLEN(instHbm_AXI_27_ARLEN),
    .AXI_27_ARSIZE(instHbm_AXI_27_ARSIZE),
    .AXI_27_ARVALID(instHbm_AXI_27_ARVALID),
    .AXI_27_ARREADY(instHbm_AXI_27_ARREADY),
    .AXI_27_AWADDR(instHbm_AXI_27_AWADDR),
    .AXI_27_AWBURST(instHbm_AXI_27_AWBURST),
    .AXI_27_AWID(instHbm_AXI_27_AWID),
    .AXI_27_AWLEN(instHbm_AXI_27_AWLEN),
    .AXI_27_AWSIZE(instHbm_AXI_27_AWSIZE),
    .AXI_27_AWVALID(instHbm_AXI_27_AWVALID),
    .AXI_27_AWREADY(instHbm_AXI_27_AWREADY),
    .AXI_27_WDATA(instHbm_AXI_27_WDATA),
    .AXI_27_WLAST(instHbm_AXI_27_WLAST),
    .AXI_27_WSTRB(instHbm_AXI_27_WSTRB),
    .AXI_27_WVALID(instHbm_AXI_27_WVALID),
    .AXI_27_WREADY(instHbm_AXI_27_WREADY),
    .AXI_27_RDATA(instHbm_AXI_27_RDATA),
    .AXI_27_RID(instHbm_AXI_27_RID),
    .AXI_27_RLAST(instHbm_AXI_27_RLAST),
    .AXI_27_RRESP(instHbm_AXI_27_RRESP),
    .AXI_27_RVALID(instHbm_AXI_27_RVALID),
    .AXI_27_RREADY(instHbm_AXI_27_RREADY),
    .AXI_27_BID(instHbm_AXI_27_BID),
    .AXI_27_BRESP(instHbm_AXI_27_BRESP),
    .AXI_27_BVALID(instHbm_AXI_27_BVALID),
    .AXI_27_BREADY(instHbm_AXI_27_BREADY),
    .AXI_27_WDATA_PARITY(instHbm_AXI_27_WDATA_PARITY),
    .AXI_27_RDATA_PARITY(instHbm_AXI_27_RDATA_PARITY),
    .AXI_28_ACLK(instHbm_AXI_28_ACLK),
    .AXI_28_ARESET_N(instHbm_AXI_28_ARESET_N),
    .AXI_28_ARADDR(instHbm_AXI_28_ARADDR),
    .AXI_28_ARBURST(instHbm_AXI_28_ARBURST),
    .AXI_28_ARID(instHbm_AXI_28_ARID),
    .AXI_28_ARLEN(instHbm_AXI_28_ARLEN),
    .AXI_28_ARSIZE(instHbm_AXI_28_ARSIZE),
    .AXI_28_ARVALID(instHbm_AXI_28_ARVALID),
    .AXI_28_ARREADY(instHbm_AXI_28_ARREADY),
    .AXI_28_AWADDR(instHbm_AXI_28_AWADDR),
    .AXI_28_AWBURST(instHbm_AXI_28_AWBURST),
    .AXI_28_AWID(instHbm_AXI_28_AWID),
    .AXI_28_AWLEN(instHbm_AXI_28_AWLEN),
    .AXI_28_AWSIZE(instHbm_AXI_28_AWSIZE),
    .AXI_28_AWVALID(instHbm_AXI_28_AWVALID),
    .AXI_28_AWREADY(instHbm_AXI_28_AWREADY),
    .AXI_28_WDATA(instHbm_AXI_28_WDATA),
    .AXI_28_WLAST(instHbm_AXI_28_WLAST),
    .AXI_28_WSTRB(instHbm_AXI_28_WSTRB),
    .AXI_28_WVALID(instHbm_AXI_28_WVALID),
    .AXI_28_WREADY(instHbm_AXI_28_WREADY),
    .AXI_28_RDATA(instHbm_AXI_28_RDATA),
    .AXI_28_RID(instHbm_AXI_28_RID),
    .AXI_28_RLAST(instHbm_AXI_28_RLAST),
    .AXI_28_RRESP(instHbm_AXI_28_RRESP),
    .AXI_28_RVALID(instHbm_AXI_28_RVALID),
    .AXI_28_RREADY(instHbm_AXI_28_RREADY),
    .AXI_28_BID(instHbm_AXI_28_BID),
    .AXI_28_BRESP(instHbm_AXI_28_BRESP),
    .AXI_28_BVALID(instHbm_AXI_28_BVALID),
    .AXI_28_BREADY(instHbm_AXI_28_BREADY),
    .AXI_28_WDATA_PARITY(instHbm_AXI_28_WDATA_PARITY),
    .AXI_28_RDATA_PARITY(instHbm_AXI_28_RDATA_PARITY),
    .AXI_29_ACLK(instHbm_AXI_29_ACLK),
    .AXI_29_ARESET_N(instHbm_AXI_29_ARESET_N),
    .AXI_29_ARADDR(instHbm_AXI_29_ARADDR),
    .AXI_29_ARBURST(instHbm_AXI_29_ARBURST),
    .AXI_29_ARID(instHbm_AXI_29_ARID),
    .AXI_29_ARLEN(instHbm_AXI_29_ARLEN),
    .AXI_29_ARSIZE(instHbm_AXI_29_ARSIZE),
    .AXI_29_ARVALID(instHbm_AXI_29_ARVALID),
    .AXI_29_ARREADY(instHbm_AXI_29_ARREADY),
    .AXI_29_AWADDR(instHbm_AXI_29_AWADDR),
    .AXI_29_AWBURST(instHbm_AXI_29_AWBURST),
    .AXI_29_AWID(instHbm_AXI_29_AWID),
    .AXI_29_AWLEN(instHbm_AXI_29_AWLEN),
    .AXI_29_AWSIZE(instHbm_AXI_29_AWSIZE),
    .AXI_29_AWVALID(instHbm_AXI_29_AWVALID),
    .AXI_29_AWREADY(instHbm_AXI_29_AWREADY),
    .AXI_29_WDATA(instHbm_AXI_29_WDATA),
    .AXI_29_WLAST(instHbm_AXI_29_WLAST),
    .AXI_29_WSTRB(instHbm_AXI_29_WSTRB),
    .AXI_29_WVALID(instHbm_AXI_29_WVALID),
    .AXI_29_WREADY(instHbm_AXI_29_WREADY),
    .AXI_29_RDATA(instHbm_AXI_29_RDATA),
    .AXI_29_RID(instHbm_AXI_29_RID),
    .AXI_29_RLAST(instHbm_AXI_29_RLAST),
    .AXI_29_RRESP(instHbm_AXI_29_RRESP),
    .AXI_29_RVALID(instHbm_AXI_29_RVALID),
    .AXI_29_RREADY(instHbm_AXI_29_RREADY),
    .AXI_29_BID(instHbm_AXI_29_BID),
    .AXI_29_BRESP(instHbm_AXI_29_BRESP),
    .AXI_29_BVALID(instHbm_AXI_29_BVALID),
    .AXI_29_BREADY(instHbm_AXI_29_BREADY),
    .AXI_29_WDATA_PARITY(instHbm_AXI_29_WDATA_PARITY),
    .AXI_29_RDATA_PARITY(instHbm_AXI_29_RDATA_PARITY),
    .AXI_30_ACLK(instHbm_AXI_30_ACLK),
    .AXI_30_ARESET_N(instHbm_AXI_30_ARESET_N),
    .AXI_30_ARADDR(instHbm_AXI_30_ARADDR),
    .AXI_30_ARBURST(instHbm_AXI_30_ARBURST),
    .AXI_30_ARID(instHbm_AXI_30_ARID),
    .AXI_30_ARLEN(instHbm_AXI_30_ARLEN),
    .AXI_30_ARSIZE(instHbm_AXI_30_ARSIZE),
    .AXI_30_ARVALID(instHbm_AXI_30_ARVALID),
    .AXI_30_ARREADY(instHbm_AXI_30_ARREADY),
    .AXI_30_AWADDR(instHbm_AXI_30_AWADDR),
    .AXI_30_AWBURST(instHbm_AXI_30_AWBURST),
    .AXI_30_AWID(instHbm_AXI_30_AWID),
    .AXI_30_AWLEN(instHbm_AXI_30_AWLEN),
    .AXI_30_AWSIZE(instHbm_AXI_30_AWSIZE),
    .AXI_30_AWVALID(instHbm_AXI_30_AWVALID),
    .AXI_30_AWREADY(instHbm_AXI_30_AWREADY),
    .AXI_30_WDATA(instHbm_AXI_30_WDATA),
    .AXI_30_WLAST(instHbm_AXI_30_WLAST),
    .AXI_30_WSTRB(instHbm_AXI_30_WSTRB),
    .AXI_30_WVALID(instHbm_AXI_30_WVALID),
    .AXI_30_WREADY(instHbm_AXI_30_WREADY),
    .AXI_30_RDATA(instHbm_AXI_30_RDATA),
    .AXI_30_RID(instHbm_AXI_30_RID),
    .AXI_30_RLAST(instHbm_AXI_30_RLAST),
    .AXI_30_RRESP(instHbm_AXI_30_RRESP),
    .AXI_30_RVALID(instHbm_AXI_30_RVALID),
    .AXI_30_RREADY(instHbm_AXI_30_RREADY),
    .AXI_30_BID(instHbm_AXI_30_BID),
    .AXI_30_BRESP(instHbm_AXI_30_BRESP),
    .AXI_30_BVALID(instHbm_AXI_30_BVALID),
    .AXI_30_BREADY(instHbm_AXI_30_BREADY),
    .AXI_30_WDATA_PARITY(instHbm_AXI_30_WDATA_PARITY),
    .AXI_30_RDATA_PARITY(instHbm_AXI_30_RDATA_PARITY),
    .AXI_31_ACLK(instHbm_AXI_31_ACLK),
    .AXI_31_ARESET_N(instHbm_AXI_31_ARESET_N),
    .AXI_31_ARADDR(instHbm_AXI_31_ARADDR),
    .AXI_31_ARBURST(instHbm_AXI_31_ARBURST),
    .AXI_31_ARID(instHbm_AXI_31_ARID),
    .AXI_31_ARLEN(instHbm_AXI_31_ARLEN),
    .AXI_31_ARSIZE(instHbm_AXI_31_ARSIZE),
    .AXI_31_ARVALID(instHbm_AXI_31_ARVALID),
    .AXI_31_ARREADY(instHbm_AXI_31_ARREADY),
    .AXI_31_AWADDR(instHbm_AXI_31_AWADDR),
    .AXI_31_AWBURST(instHbm_AXI_31_AWBURST),
    .AXI_31_AWID(instHbm_AXI_31_AWID),
    .AXI_31_AWLEN(instHbm_AXI_31_AWLEN),
    .AXI_31_AWSIZE(instHbm_AXI_31_AWSIZE),
    .AXI_31_AWVALID(instHbm_AXI_31_AWVALID),
    .AXI_31_AWREADY(instHbm_AXI_31_AWREADY),
    .AXI_31_WDATA(instHbm_AXI_31_WDATA),
    .AXI_31_WLAST(instHbm_AXI_31_WLAST),
    .AXI_31_WSTRB(instHbm_AXI_31_WSTRB),
    .AXI_31_WVALID(instHbm_AXI_31_WVALID),
    .AXI_31_WREADY(instHbm_AXI_31_WREADY),
    .AXI_31_RDATA(instHbm_AXI_31_RDATA),
    .AXI_31_RID(instHbm_AXI_31_RID),
    .AXI_31_RLAST(instHbm_AXI_31_RLAST),
    .AXI_31_RRESP(instHbm_AXI_31_RRESP),
    .AXI_31_RVALID(instHbm_AXI_31_RVALID),
    .AXI_31_RREADY(instHbm_AXI_31_RREADY),
    .AXI_31_BID(instHbm_AXI_31_BID),
    .AXI_31_BRESP(instHbm_AXI_31_BRESP),
    .AXI_31_BVALID(instHbm_AXI_31_BVALID),
    .AXI_31_BREADY(instHbm_AXI_31_BREADY),
    .AXI_31_WDATA_PARITY(instHbm_AXI_31_WDATA_PARITY),
    .AXI_31_RDATA_PARITY(instHbm_AXI_31_RDATA_PARITY),
    .APB_0_PWDATA(instHbm_APB_0_PWDATA),
    .APB_0_PADDR(instHbm_APB_0_PADDR),
    .APB_0_PCLK(instHbm_APB_0_PCLK),
    .APB_0_PENABLE(instHbm_APB_0_PENABLE),
    .APB_0_PRESET_N(instHbm_APB_0_PRESET_N),
    .APB_0_PSEL(instHbm_APB_0_PSEL),
    .APB_0_PWRITE(instHbm_APB_0_PWRITE),
    .APB_0_PRDATA(instHbm_APB_0_PRDATA),
    .APB_0_PREADY(instHbm_APB_0_PREADY),
    .APB_0_PSLVERR(instHbm_APB_0_PSLVERR),
    .APB_1_PWDATA(instHbm_APB_1_PWDATA),
    .APB_1_PADDR(instHbm_APB_1_PADDR),
    .APB_1_PCLK(instHbm_APB_1_PCLK),
    .APB_1_PENABLE(instHbm_APB_1_PENABLE),
    .APB_1_PRESET_N(instHbm_APB_1_PRESET_N),
    .APB_1_PSEL(instHbm_APB_1_PSEL),
    .APB_1_PWRITE(instHbm_APB_1_PWRITE),
    .APB_1_PRDATA(instHbm_APB_1_PRDATA),
    .APB_1_PREADY(instHbm_APB_1_PREADY),
    .APB_1_PSLVERR(instHbm_APB_1_PSLVERR),
    .DRAM_0_STAT_CATTRIP(instHbm_DRAM_0_STAT_CATTRIP),
    .DRAM_0_STAT_TEMP(instHbm_DRAM_0_STAT_TEMP),
    .DRAM_1_STAT_CATTRIP(instHbm_DRAM_1_STAT_CATTRIP),
    .DRAM_1_STAT_TEMP(instHbm_DRAM_1_STAT_TEMP),
    .apb_complete_0(instHbm_apb_complete_0),
    .apb_complete_1(instHbm_apb_complete_1)
  );
  assign io_hbm_clk = axiAclk_pad_O; // @[HBMDriver.scala 90:25]
  assign io_hbm_rstn = _io_hbm_rstn_T_2 & apb_complete_1; // @[HBMDriver.scala 99:17]
  assign io_axi_hbm_0_aw_ready = instHbm_AXI_00_AWREADY; // @[HBMDriver.scala 32:32 HBMDriver.scala 130:49]
  assign io_axi_hbm_0_ar_ready = instHbm_AXI_00_ARREADY; // @[HBMDriver.scala 32:32 HBMDriver.scala 123:49]
  assign io_axi_hbm_0_w_ready = instHbm_AXI_00_WREADY; // @[HBMDriver.scala 32:32 HBMDriver.scala 135:49]
  assign io_axi_hbm_0_r_valid = instHbm_AXI_00_RVALID; // @[HBMDriver.scala 32:32 HBMDriver.scala 140:49]
  assign io_axi_hbm_0_r_bits_data = instHbm_AXI_00_RDATA; // @[HBMDriver.scala 32:32 HBMDriver.scala 136:49]
  assign io_axi_hbm_1_aw_ready = instHbm_AXI_01_AWREADY; // @[HBMDriver.scala 32:32 HBMDriver.scala 164:49]
  assign io_axi_hbm_1_ar_ready = instHbm_AXI_01_ARREADY; // @[HBMDriver.scala 32:32 HBMDriver.scala 157:49]
  assign io_axi_hbm_1_w_ready = instHbm_AXI_01_WREADY; // @[HBMDriver.scala 32:32 HBMDriver.scala 169:49]
  assign io_axi_hbm_1_r_valid = instHbm_AXI_01_RVALID; // @[HBMDriver.scala 32:32 HBMDriver.scala 174:49]
  assign io_axi_hbm_1_r_bits_data = instHbm_AXI_01_RDATA; // @[HBMDriver.scala 32:32 HBMDriver.scala 170:49]
  assign io_axi_hbm_1_r_bits_last = instHbm_AXI_01_RLAST; // @[HBMDriver.scala 32:32 HBMDriver.scala 172:49]
  assign io_axi_hbm_1_b_valid = instHbm_AXI_01_BVALID; // @[HBMDriver.scala 32:32 HBMDriver.scala 178:49]
  assign mmcmGlbl_io_CLKIN1 = clock; // @[HBMDriver.scala 60:33]
  assign apb0Pclk_pad_I = mmcmGlbl_io_CLKOUT0; // @[Buf.scala 34:26]
  assign apb0Pclk_pad_1_I = apb0Pclk_pad_O; // @[HBMDriver.scala 63:63]
  assign apb0Pclk_pad_2_I = apb0Pclk_pad_1_O; // @[HBMDriver.scala 63:71]
  assign axiAclkIn0_pad_I = mmcmGlbl_io_CLKOUT1; // @[Buf.scala 34:26]
  assign hbmRefClk0_pad_I = mmcmGlbl_io_CLKOUT2; // @[Buf.scala 34:26]
  assign apb1Pclk_pad_I = mmcmGlbl_io_CLKOUT3; // @[Buf.scala 34:26]
  assign apb1Pclk_pad_1_I = apb1Pclk_pad_O; // @[HBMDriver.scala 66:63]
  assign apb1Pclk_pad_2_I = apb1Pclk_pad_1_O; // @[HBMDriver.scala 66:71]
  assign axiAclkIn1_pad_I = mmcmGlbl_io_CLKOUT4; // @[Buf.scala 34:26]
  assign hbmRefClk1_pad_I = mmcmGlbl_io_CLKOUT5; // @[Buf.scala 34:26]
  assign mmcmAxi_io_CLKIN1 = axiAclkIn0_pad_O; // @[HBMDriver.scala 84:33]
  assign mmcmAxi_io_RST = ~mmcmGlbl_io_LOCKED; // @[HBMDriver.scala 85:36]
  assign axiAclk_pad_I = mmcmAxi_io_CLKOUT0; // @[Buf.scala 34:26]
  assign instHbm_HBM_REF_CLK_0 = hbmRefClk0_pad_O; // @[HBMDriver.scala 103:41]
  assign instHbm_HBM_REF_CLK_1 = hbmRefClk1_pad_O; // @[HBMDriver.scala 104:41]
  assign instHbm_AXI_00_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 115:49]
  assign instHbm_AXI_00_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 116:49]
  assign instHbm_AXI_00_ARADDR = io_axi_hbm_0_ar_bits_addr[32:0]; // @[HBMDriver.scala 117:49]
  assign instHbm_AXI_00_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARLEN = io_axi_hbm_0_ar_bits_len; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_ARVALID = io_axi_hbm_0_ar_valid; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWADDR = io_axi_hbm_0_aw_bits_addr[32:0]; // @[HBMDriver.scala 124:49]
  assign instHbm_AXI_00_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWLEN = io_axi_hbm_0_aw_bits_len; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_AWVALID = io_axi_hbm_0_aw_valid; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WDATA = io_axi_hbm_0_w_bits_data; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WLAST = io_axi_hbm_0_w_bits_last; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WVALID = io_axi_hbm_0_w_valid; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_RREADY = io_axi_hbm_0_r_ready; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_00_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 146:49]
  assign instHbm_AXI_01_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 149:49]
  assign instHbm_AXI_01_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 150:49]
  assign instHbm_AXI_01_ARADDR = io_axi_hbm_1_ar_bits_addr[32:0]; // @[HBMDriver.scala 151:49]
  assign instHbm_AXI_01_ARBURST = io_axi_hbm_1_ar_bits_burst; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARLEN = io_axi_hbm_1_ar_bits_len; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARSIZE = io_axi_hbm_1_ar_bits_size; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_ARVALID = io_axi_hbm_1_ar_valid; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWADDR = io_axi_hbm_1_aw_bits_addr[32:0]; // @[HBMDriver.scala 158:49]
  assign instHbm_AXI_01_AWBURST = io_axi_hbm_1_aw_bits_burst; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWLEN = io_axi_hbm_1_aw_bits_len; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWSIZE = io_axi_hbm_1_aw_bits_size; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_AWVALID = io_axi_hbm_1_aw_valid; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WDATA = io_axi_hbm_1_w_bits_data; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WLAST = io_axi_hbm_1_w_bits_last; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WSTRB = io_axi_hbm_1_w_bits_strb; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WVALID = io_axi_hbm_1_w_valid; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_RREADY = io_axi_hbm_1_r_ready; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_BREADY = io_axi_hbm_1_b_ready; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_01_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 180:49]
  assign instHbm_AXI_02_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 183:49]
  assign instHbm_AXI_02_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 184:49]
  assign instHbm_AXI_02_ARADDR = 33'h0; // @[HBMDriver.scala 185:49]
  assign instHbm_AXI_02_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWADDR = 33'h0; // @[HBMDriver.scala 192:49]
  assign instHbm_AXI_02_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_02_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 214:49]
  assign instHbm_AXI_03_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 217:49]
  assign instHbm_AXI_03_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 218:49]
  assign instHbm_AXI_03_ARADDR = 33'h0; // @[HBMDriver.scala 219:49]
  assign instHbm_AXI_03_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWADDR = 33'h0; // @[HBMDriver.scala 226:49]
  assign instHbm_AXI_03_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_03_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 248:49]
  assign instHbm_AXI_04_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 251:49]
  assign instHbm_AXI_04_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 252:49]
  assign instHbm_AXI_04_ARADDR = 33'h0; // @[HBMDriver.scala 253:49]
  assign instHbm_AXI_04_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWADDR = 33'h0; // @[HBMDriver.scala 260:49]
  assign instHbm_AXI_04_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_04_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 282:49]
  assign instHbm_AXI_05_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 285:49]
  assign instHbm_AXI_05_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 286:49]
  assign instHbm_AXI_05_ARADDR = 33'h0; // @[HBMDriver.scala 287:49]
  assign instHbm_AXI_05_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWADDR = 33'h0; // @[HBMDriver.scala 294:49]
  assign instHbm_AXI_05_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_05_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 316:49]
  assign instHbm_AXI_06_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 319:49]
  assign instHbm_AXI_06_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 320:49]
  assign instHbm_AXI_06_ARADDR = 33'h0; // @[HBMDriver.scala 321:49]
  assign instHbm_AXI_06_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWADDR = 33'h0; // @[HBMDriver.scala 328:49]
  assign instHbm_AXI_06_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_06_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 350:49]
  assign instHbm_AXI_07_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 353:49]
  assign instHbm_AXI_07_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 354:49]
  assign instHbm_AXI_07_ARADDR = 33'h0; // @[HBMDriver.scala 355:49]
  assign instHbm_AXI_07_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWADDR = 33'h0; // @[HBMDriver.scala 362:49]
  assign instHbm_AXI_07_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_07_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 384:49]
  assign instHbm_AXI_08_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 387:49]
  assign instHbm_AXI_08_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 388:49]
  assign instHbm_AXI_08_ARADDR = 33'h0; // @[HBMDriver.scala 389:49]
  assign instHbm_AXI_08_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWADDR = 33'h0; // @[HBMDriver.scala 396:49]
  assign instHbm_AXI_08_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_08_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 418:49]
  assign instHbm_AXI_09_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 421:49]
  assign instHbm_AXI_09_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 422:49]
  assign instHbm_AXI_09_ARADDR = 33'h0; // @[HBMDriver.scala 423:49]
  assign instHbm_AXI_09_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWADDR = 33'h0; // @[HBMDriver.scala 430:49]
  assign instHbm_AXI_09_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_09_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 452:49]
  assign instHbm_AXI_10_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 455:49]
  assign instHbm_AXI_10_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 456:49]
  assign instHbm_AXI_10_ARADDR = 33'h0; // @[HBMDriver.scala 457:49]
  assign instHbm_AXI_10_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWADDR = 33'h0; // @[HBMDriver.scala 464:49]
  assign instHbm_AXI_10_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_10_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 486:49]
  assign instHbm_AXI_11_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 489:49]
  assign instHbm_AXI_11_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 490:49]
  assign instHbm_AXI_11_ARADDR = 33'h0; // @[HBMDriver.scala 491:49]
  assign instHbm_AXI_11_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWADDR = 33'h0; // @[HBMDriver.scala 498:49]
  assign instHbm_AXI_11_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_11_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 520:49]
  assign instHbm_AXI_12_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 523:49]
  assign instHbm_AXI_12_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 524:49]
  assign instHbm_AXI_12_ARADDR = 33'h0; // @[HBMDriver.scala 525:49]
  assign instHbm_AXI_12_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWADDR = 33'h0; // @[HBMDriver.scala 532:49]
  assign instHbm_AXI_12_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_12_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 554:49]
  assign instHbm_AXI_13_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 557:49]
  assign instHbm_AXI_13_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 558:49]
  assign instHbm_AXI_13_ARADDR = 33'h0; // @[HBMDriver.scala 559:49]
  assign instHbm_AXI_13_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWADDR = 33'h0; // @[HBMDriver.scala 566:49]
  assign instHbm_AXI_13_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_13_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 588:49]
  assign instHbm_AXI_14_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 591:49]
  assign instHbm_AXI_14_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 592:49]
  assign instHbm_AXI_14_ARADDR = 33'h0; // @[HBMDriver.scala 593:49]
  assign instHbm_AXI_14_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWADDR = 33'h0; // @[HBMDriver.scala 600:49]
  assign instHbm_AXI_14_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_14_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 622:49]
  assign instHbm_AXI_15_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 625:49]
  assign instHbm_AXI_15_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 626:49]
  assign instHbm_AXI_15_ARADDR = 33'h0; // @[HBMDriver.scala 627:49]
  assign instHbm_AXI_15_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWADDR = 33'h0; // @[HBMDriver.scala 634:49]
  assign instHbm_AXI_15_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_15_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 656:49]
  assign instHbm_AXI_16_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 667:49]
  assign instHbm_AXI_16_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 668:49]
  assign instHbm_AXI_16_ARADDR = 33'h0; // @[HBMDriver.scala 669:49]
  assign instHbm_AXI_16_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWADDR = 33'h0; // @[HBMDriver.scala 676:49]
  assign instHbm_AXI_16_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_16_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 698:49]
  assign instHbm_AXI_17_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 701:49]
  assign instHbm_AXI_17_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 702:49]
  assign instHbm_AXI_17_ARADDR = 33'h0; // @[HBMDriver.scala 703:49]
  assign instHbm_AXI_17_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWADDR = 33'h0; // @[HBMDriver.scala 710:49]
  assign instHbm_AXI_17_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_17_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 732:49]
  assign instHbm_AXI_18_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 735:49]
  assign instHbm_AXI_18_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 736:49]
  assign instHbm_AXI_18_ARADDR = 33'h0; // @[HBMDriver.scala 737:49]
  assign instHbm_AXI_18_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWADDR = 33'h0; // @[HBMDriver.scala 744:49]
  assign instHbm_AXI_18_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_18_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 766:49]
  assign instHbm_AXI_19_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 769:49]
  assign instHbm_AXI_19_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 770:49]
  assign instHbm_AXI_19_ARADDR = 33'h0; // @[HBMDriver.scala 771:49]
  assign instHbm_AXI_19_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWADDR = 33'h0; // @[HBMDriver.scala 778:49]
  assign instHbm_AXI_19_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_19_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 800:49]
  assign instHbm_AXI_20_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 803:49]
  assign instHbm_AXI_20_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 804:49]
  assign instHbm_AXI_20_ARADDR = 33'h0; // @[HBMDriver.scala 805:49]
  assign instHbm_AXI_20_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWADDR = 33'h0; // @[HBMDriver.scala 812:49]
  assign instHbm_AXI_20_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_20_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 834:49]
  assign instHbm_AXI_21_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 837:49]
  assign instHbm_AXI_21_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 838:49]
  assign instHbm_AXI_21_ARADDR = 33'h0; // @[HBMDriver.scala 839:49]
  assign instHbm_AXI_21_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWADDR = 33'h0; // @[HBMDriver.scala 846:49]
  assign instHbm_AXI_21_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_21_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 868:49]
  assign instHbm_AXI_22_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 871:49]
  assign instHbm_AXI_22_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 872:49]
  assign instHbm_AXI_22_ARADDR = 33'h0; // @[HBMDriver.scala 873:49]
  assign instHbm_AXI_22_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWADDR = 33'h0; // @[HBMDriver.scala 880:49]
  assign instHbm_AXI_22_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_22_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 902:49]
  assign instHbm_AXI_23_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 905:49]
  assign instHbm_AXI_23_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 906:49]
  assign instHbm_AXI_23_ARADDR = 33'h0; // @[HBMDriver.scala 907:49]
  assign instHbm_AXI_23_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWADDR = 33'h0; // @[HBMDriver.scala 914:49]
  assign instHbm_AXI_23_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_23_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 936:49]
  assign instHbm_AXI_24_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 939:49]
  assign instHbm_AXI_24_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 940:49]
  assign instHbm_AXI_24_ARADDR = 33'h0; // @[HBMDriver.scala 941:49]
  assign instHbm_AXI_24_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWADDR = 33'h0; // @[HBMDriver.scala 948:49]
  assign instHbm_AXI_24_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_24_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 970:49]
  assign instHbm_AXI_25_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 973:49]
  assign instHbm_AXI_25_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 974:49]
  assign instHbm_AXI_25_ARADDR = 33'h0; // @[HBMDriver.scala 975:49]
  assign instHbm_AXI_25_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWADDR = 33'h0; // @[HBMDriver.scala 982:49]
  assign instHbm_AXI_25_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_25_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1004:49]
  assign instHbm_AXI_26_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1007:49]
  assign instHbm_AXI_26_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1008:49]
  assign instHbm_AXI_26_ARADDR = 33'h0; // @[HBMDriver.scala 1009:49]
  assign instHbm_AXI_26_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWADDR = 33'h0; // @[HBMDriver.scala 1016:49]
  assign instHbm_AXI_26_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_26_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1038:49]
  assign instHbm_AXI_27_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1041:49]
  assign instHbm_AXI_27_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1042:49]
  assign instHbm_AXI_27_ARADDR = 33'h0; // @[HBMDriver.scala 1043:49]
  assign instHbm_AXI_27_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWADDR = 33'h0; // @[HBMDriver.scala 1050:49]
  assign instHbm_AXI_27_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_27_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1072:49]
  assign instHbm_AXI_28_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1075:49]
  assign instHbm_AXI_28_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1076:49]
  assign instHbm_AXI_28_ARADDR = 33'h0; // @[HBMDriver.scala 1077:49]
  assign instHbm_AXI_28_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWADDR = 33'h0; // @[HBMDriver.scala 1084:49]
  assign instHbm_AXI_28_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_28_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1106:49]
  assign instHbm_AXI_29_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1109:49]
  assign instHbm_AXI_29_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1110:49]
  assign instHbm_AXI_29_ARADDR = 33'h0; // @[HBMDriver.scala 1111:49]
  assign instHbm_AXI_29_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWADDR = 33'h0; // @[HBMDriver.scala 1118:49]
  assign instHbm_AXI_29_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_29_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1140:49]
  assign instHbm_AXI_30_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1143:49]
  assign instHbm_AXI_30_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1144:49]
  assign instHbm_AXI_30_ARADDR = 33'h0; // @[HBMDriver.scala 1145:49]
  assign instHbm_AXI_30_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWADDR = 33'h0; // @[HBMDriver.scala 1152:49]
  assign instHbm_AXI_30_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_30_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1174:49]
  assign instHbm_AXI_31_ACLK = axiAclk_pad_O; // @[HBMDriver.scala 1177:49]
  assign instHbm_AXI_31_ARESET_N = mmcmAxi_io_LOCKED; // @[HBMDriver.scala 1178:49]
  assign instHbm_AXI_31_ARADDR = 33'h0; // @[HBMDriver.scala 1179:49]
  assign instHbm_AXI_31_ARBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_ARVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWADDR = 33'h0; // @[HBMDriver.scala 1186:49]
  assign instHbm_AXI_31_AWBURST = 2'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWID = 6'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWLEN = 4'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWSIZE = 3'h5; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_AWVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WDATA = 256'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WLAST = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WSTRB = 32'hffffffff; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WVALID = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_RREADY = 1'h0; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_BREADY = 1'h1; // @[HBMDriver.scala 32:32 HBMDriver.scala 42:39]
  assign instHbm_AXI_31_WDATA_PARITY = 32'h0; // @[HBMDriver.scala 1208:49]
  assign instHbm_APB_0_PWDATA = 32'h0; // @[HBMDriver.scala 1214:36]
  assign instHbm_APB_0_PADDR = 22'h0; // @[HBMDriver.scala 1215:36]
  assign instHbm_APB_0_PCLK = apb0Pclk_pad_2_O; // @[HBMDriver.scala 1216:36]
  assign instHbm_APB_0_PENABLE = 1'h0; // @[HBMDriver.scala 1217:36]
  assign instHbm_APB_0_PRESET_N = mmcmGlbl_io_LOCKED; // @[HBMDriver.scala 1218:36]
  assign instHbm_APB_0_PSEL = 1'h0; // @[HBMDriver.scala 1219:36]
  assign instHbm_APB_0_PWRITE = 1'h0; // @[HBMDriver.scala 1220:36]
  assign instHbm_APB_1_PWDATA = 32'h0; // @[HBMDriver.scala 1225:36]
  assign instHbm_APB_1_PADDR = 22'h0; // @[HBMDriver.scala 1226:36]
  assign instHbm_APB_1_PCLK = apb1Pclk_pad_2_O; // @[HBMDriver.scala 1227:36]
  assign instHbm_APB_1_PENABLE = 1'h0; // @[HBMDriver.scala 1228:36]
  assign instHbm_APB_1_PRESET_N = mmcmGlbl_io_LOCKED; // @[HBMDriver.scala 1229:36]
  assign instHbm_APB_1_PSEL = 1'h0; // @[HBMDriver.scala 1230:36]
  assign instHbm_APB_1_PWRITE = 1'h0; // @[HBMDriver.scala 1231:36]
  always @(posedge apb0Pclk_pad_2_O) begin
    apb_complete_0_r <= instHbm_apb_complete_0; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    apb_complete_0 <= apb_complete_0_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  end
  always @(posedge apb1Pclk_pad_2_O) begin
    apb_complete_1_r <= instHbm_apb_complete_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    apb_complete_1 <= apb_complete_1_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  end
  always @(posedge axiAclk_pad_O) begin
    io_hbm_rstn_REG <= mmcmAxi_io_LOCKED; // @[HBMDriver.scala 97:63]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  apb_complete_0_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  apb_complete_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  apb_complete_1_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  apb_complete_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_hbm_rstn_REG = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SV_STREAM_FIFO(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [599:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [599:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [599:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [74:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [599:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [74:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [74:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(600), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 75'h7ffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 75'h7ffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter(
  input          io_in_clk,
  input          io_out_clk,
  input          io_rstn,
  output         io_in_ready,
  input          io_in_valid,
  input  [511:0] io_in_bits_data,
  input  [31:0]  io_in_bits_tcrc,
  input  [10:0]  io_in_bits_tuser_qid,
  input  [2:0]   io_in_bits_tuser_port_id,
  input          io_in_bits_tuser_err,
  input  [31:0]  io_in_bits_tuser_mdata,
  input  [5:0]   io_in_bits_tuser_mty,
  input          io_in_bits_tuser_zero_byte,
  input          io_in_bits_last,
  input          io_out_ready,
  output         io_out_valid,
  output [511:0] io_out_bits_data
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [599:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [599:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [598:0] _fifo_io_in_data_T = {io_in_bits_data,io_in_bits_tcrc,io_in_bits_tuser_qid,io_in_bits_tuser_port_id,
    io_in_bits_tuser_err,io_in_bits_tuser_mdata,io_in_bits_tuser_mty,io_in_bits_tuser_zero_byte,io_in_bits_last}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_data = fifo_io_out_data[598:87]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{1'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module SV_STREAM_FIFO_1(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [607:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [607:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [607:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [75:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [607:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [75:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [75:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(608), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 76'hfffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 76'hfffffffffffffffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_1(
  input          io_in_clk,
  input          io_out_clk,
  input          io_rstn,
  output         io_in_ready,
  input          io_in_valid,
  input  [511:0] io_in_bits_data,
  input  [31:0]  io_in_bits_tcrc,
  input          io_in_bits_ctrl_marker,
  input  [6:0]   io_in_bits_ctrl_ecc,
  input  [31:0]  io_in_bits_ctrl_len,
  input  [2:0]   io_in_bits_ctrl_port_id,
  input  [10:0]  io_in_bits_ctrl_qid,
  input          io_in_bits_ctrl_has_cmpt,
  input          io_in_bits_last,
  input  [5:0]   io_in_bits_mty,
  input          io_out_ready,
  output         io_out_valid,
  output [511:0] io_out_bits_data,
  output [31:0]  io_out_bits_tcrc,
  output         io_out_bits_ctrl_marker,
  output [6:0]   io_out_bits_ctrl_ecc,
  output [31:0]  io_out_bits_ctrl_len,
  output [2:0]   io_out_bits_ctrl_port_id,
  output [10:0]  io_out_bits_ctrl_qid,
  output         io_out_bits_ctrl_has_cmpt,
  output         io_out_bits_last,
  output [5:0]   io_out_bits_mty
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [607:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [607:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [605:0] _fifo_io_in_data_T = {io_in_bits_data,io_in_bits_tcrc,io_in_bits_ctrl_marker,io_in_bits_ctrl_ecc,
    io_in_bits_ctrl_len,io_in_bits_ctrl_port_id,io_in_bits_ctrl_qid,io_in_bits_ctrl_has_cmpt,io_in_bits_last,
    io_in_bits_mty}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_1 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_data = fifo_io_out_data[605:94]; // @[XConverter.scala 107:77]
  assign io_out_bits_tcrc = fifo_io_out_data[93:62]; // @[XConverter.scala 107:77]
  assign io_out_bits_ctrl_marker = fifo_io_out_data[61]; // @[XConverter.scala 107:77]
  assign io_out_bits_ctrl_ecc = fifo_io_out_data[60:54]; // @[XConverter.scala 107:77]
  assign io_out_bits_ctrl_len = fifo_io_out_data[53:22]; // @[XConverter.scala 107:77]
  assign io_out_bits_ctrl_port_id = fifo_io_out_data[21:19]; // @[XConverter.scala 107:77]
  assign io_out_bits_ctrl_qid = fifo_io_out_data[18:8]; // @[XConverter.scala 107:77]
  assign io_out_bits_ctrl_has_cmpt = fifo_io_out_data[7]; // @[XConverter.scala 107:77]
  assign io_out_bits_last = fifo_io_out_data[6]; // @[XConverter.scala 107:77]
  assign io_out_bits_mty = fifo_io_out_data[5:0]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{2'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module SV_STREAM_FIFO_2(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [143:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [143:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [143:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [17:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [143:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [17:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [17:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(144), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 18'h3ffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 18'h3ffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_2(
  input         io_in_clk,
  input         io_out_clk,
  input         io_rstn,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [31:0] io_in_bits_len,
  input         io_in_bits_eop,
  input         io_in_bits_sop,
  input         io_in_bits_mrkr_req,
  input         io_in_bits_sdi,
  input  [10:0] io_in_bits_qid,
  input         io_in_bits_error,
  input  [7:0]  io_in_bits_func,
  input  [15:0] io_in_bits_cidx,
  input  [2:0]  io_in_bits_port_id,
  input         io_in_bits_no_dma,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [31:0] io_out_bits_len,
  output        io_out_bits_eop,
  output        io_out_bits_sop,
  output        io_out_bits_mrkr_req,
  output        io_out_bits_sdi,
  output [10:0] io_out_bits_qid,
  output        io_out_bits_error,
  output [7:0]  io_out_bits_func,
  output [15:0] io_out_bits_cidx,
  output [2:0]  io_out_bits_port_id,
  output        io_out_bits_no_dma
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [143:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [143:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [39:0] fifo_io_in_data_lo = {io_in_bits_qid,io_in_bits_error,io_in_bits_func,io_in_bits_cidx,io_in_bits_port_id,
    io_in_bits_no_dma}; // @[XConverter.scala 103:63]
  wire [139:0] _fifo_io_in_data_T = {io_in_bits_addr,io_in_bits_len,io_in_bits_eop,io_in_bits_sop,io_in_bits_mrkr_req,
    io_in_bits_sdi,fifo_io_in_data_lo}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_2 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_addr = fifo_io_out_data[139:76]; // @[XConverter.scala 107:77]
  assign io_out_bits_len = fifo_io_out_data[75:44]; // @[XConverter.scala 107:77]
  assign io_out_bits_eop = fifo_io_out_data[43]; // @[XConverter.scala 107:77]
  assign io_out_bits_sop = fifo_io_out_data[42]; // @[XConverter.scala 107:77]
  assign io_out_bits_mrkr_req = fifo_io_out_data[41]; // @[XConverter.scala 107:77]
  assign io_out_bits_sdi = fifo_io_out_data[40]; // @[XConverter.scala 107:77]
  assign io_out_bits_qid = fifo_io_out_data[39:29]; // @[XConverter.scala 107:77]
  assign io_out_bits_error = fifo_io_out_data[28]; // @[XConverter.scala 107:77]
  assign io_out_bits_func = fifo_io_out_data[27:20]; // @[XConverter.scala 107:77]
  assign io_out_bits_cidx = fifo_io_out_data[19:4]; // @[XConverter.scala 107:77]
  assign io_out_bits_port_id = fifo_io_out_data[3:1]; // @[XConverter.scala 107:77]
  assign io_out_bits_no_dma = fifo_io_out_data[0]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{4'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module SV_STREAM_FIFO_3(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [127:0] io_in_data,
  input          io_in_valid,
  output         io_in_ready,
  output [127:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [127:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [15:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [127:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [15:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [15:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(128), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_in_ready = meta_s_axis_tready; // @[Meta.scala 34:41]
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 16'hffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 16'hffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_3(
  input         io_in_clk,
  input         io_out_clk,
  input         io_rstn,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [10:0] io_in_bits_qid,
  input         io_in_bits_error,
  input  [7:0]  io_in_bits_func,
  input  [2:0]  io_in_bits_port_id,
  input  [6:0]  io_in_bits_pfch_tag,
  input  [31:0] io_in_bits_len,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [10:0] io_out_bits_qid,
  output        io_out_bits_error,
  output [7:0]  io_out_bits_func,
  output [2:0]  io_out_bits_port_id,
  output [6:0]  io_out_bits_pfch_tag
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [127:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_in_ready; // @[XConverter.scala 97:34]
  wire [127:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire  fifo_io_out_ready; // @[XConverter.scala 97:34]
  wire [125:0] _fifo_io_in_data_T = {io_in_bits_addr,io_in_bits_qid,io_in_bits_error,io_in_bits_func,io_in_bits_port_id,
    io_in_bits_pfch_tag,io_in_bits_len}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_3 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_in_ready(fifo_io_in_ready),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_in_ready = fifo_io_in_ready; // @[XConverter.scala 105:41]
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_addr = fifo_io_out_data[125:62]; // @[XConverter.scala 107:77]
  assign io_out_bits_qid = fifo_io_out_data[61:51]; // @[XConverter.scala 107:77]
  assign io_out_bits_error = fifo_io_out_data[50]; // @[XConverter.scala 107:77]
  assign io_out_bits_func = fifo_io_out_data[49:42]; // @[XConverter.scala 107:77]
  assign io_out_bits_port_id = fifo_io_out_data[41:39]; // @[XConverter.scala 107:77]
  assign io_out_bits_pfch_tag = fifo_io_out_data[38:32]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{2'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
  assign fifo_io_out_ready = io_out_ready; // @[XConverter.scala 109:41]
endmodule
module CMDBoundaryCheck(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [6:0]  io_in_bits_pfch_tag,
  input  [31:0] io_in_bits_len,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [6:0]  io_out_bits_pfch_tag,
  output [31:0] io_out_bits_len
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [23:0] offset_addr; // @[CheckSplit.scala 129:34]
  reg [23:0] new_length; // @[CheckSplit.scala 130:33]
  reg [63:0] cmd_addr; // @[CheckSplit.scala 131:31]
  reg [31:0] cmd_len; // @[CheckSplit.scala 132:30]
  reg [63:0] mini_addr; // @[CheckSplit.scala 133:32]
  reg [31:0] mini_len; // @[CheckSplit.scala 134:31]
  reg [6:0] cmd_temp_pfch_tag; // @[CheckSplit.scala 135:27]
  reg [2:0] state; // @[CheckSplit.scala 138:28]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _offset_addr_T = io_in_bits_addr & 64'h1fffff; // @[CheckSplit.scala 154:100]
  wire [63:0] _new_length_T_2 = 64'h200000 - _offset_addr_T; // @[CheckSplit.scala 156:96]
  wire [63:0] _GEN_9 = _T_1 ? _offset_addr_T : {{40'd0}, offset_addr}; // @[CheckSplit.scala 150:43 CheckSplit.scala 154:81 CheckSplit.scala 129:34]
  wire [63:0] _GEN_11 = _T_1 ? _new_length_T_2 : {{40'd0}, new_length}; // @[CheckSplit.scala 150:43 CheckSplit.scala 156:81 CheckSplit.scala 130:33]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_143 = {{8'd0}, offset_addr}; // @[CheckSplit.scala 160:43]
  wire [31:0] _T_4 = _GEN_143 + cmd_len; // @[CheckSplit.scala 160:43]
  wire [63:0] _GEN_144 = {{40'd0}, new_length}; // @[CheckSplit.scala 163:93]
  wire [63:0] _cmd_addr_T_1 = cmd_addr + _GEN_144; // @[CheckSplit.scala 163:93]
  wire [31:0] _GEN_145 = {{8'd0}, new_length}; // @[CheckSplit.scala 164:92]
  wire [31:0] _cmd_len_T_1 = cmd_len - _GEN_145; // @[CheckSplit.scala 164:92]
  wire  _T_6 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _cmd_addr_T_3 = cmd_addr + 64'h200000; // @[CheckSplit.scala 176:93]
  wire [31:0] _cmd_len_T_3 = cmd_len - 32'h200000; // @[CheckSplit.scala 177:92]
  wire [31:0] _GEN_18 = cmd_len > 32'h200000 ? 32'h200000 : cmd_len; // @[CheckSplit.scala 173:52 CheckSplit.scala 175:81 CheckSplit.scala 181:81]
  wire [63:0] _GEN_19 = cmd_len > 32'h200000 ? _cmd_addr_T_3 : cmd_addr; // @[CheckSplit.scala 173:52 CheckSplit.scala 176:81 CheckSplit.scala 131:31]
  wire [31:0] _GEN_20 = cmd_len > 32'h200000 ? _cmd_len_T_3 : cmd_len; // @[CheckSplit.scala 173:52 CheckSplit.scala 177:81 CheckSplit.scala 132:30]
  wire [2:0] _GEN_21 = cmd_len > 32'h200000 ? 3'h3 : 3'h4; // @[CheckSplit.scala 173:52 CheckSplit.scala 178:65 CheckSplit.scala 182:65]
  wire  _T_8 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = mini_len > 32'h1000; // @[CheckSplit.scala 188:47]
  wire [63:0] _mini_addr_T_1 = mini_addr + 64'h1000; // @[CheckSplit.scala 189:94]
  wire [31:0] _mini_len_T_1 = mini_len - 32'h1000; // @[CheckSplit.scala 190:93]
  wire [63:0] _GEN_22 = mini_len > 32'h1000 ? _mini_addr_T_1 : mini_addr; // @[CheckSplit.scala 188:66 CheckSplit.scala 189:81 CheckSplit.scala 133:32]
  wire [31:0] _GEN_23 = mini_len > 32'h1000 ? _mini_len_T_1 : mini_len; // @[CheckSplit.scala 188:66 CheckSplit.scala 190:81 CheckSplit.scala 134:31]
  wire [31:0] _GEN_25 = mini_len > 32'h1000 ? 32'h1000 : mini_len; // @[CheckSplit.scala 188:66 CheckSplit.scala 193:73 CheckSplit.scala 198:73]
  wire [2:0] _GEN_32 = mini_len > 32'h1000 ? state : 3'h2; // @[CheckSplit.scala 188:66 CheckSplit.scala 138:28 CheckSplit.scala 200:81]
  wire [63:0] _GEN_34 = io_out_ready ? _GEN_22 : mini_addr; // @[CheckSplit.scala 186:51 CheckSplit.scala 133:32]
  wire [31:0] _GEN_35 = io_out_ready ? _GEN_23 : mini_len; // @[CheckSplit.scala 186:51 CheckSplit.scala 134:31]
  wire [31:0] _GEN_37 = io_out_ready ? _GEN_25 : 32'h0; // @[CheckSplit.scala 186:51 CheckSplit.scala 143:33]
  wire [6:0] _GEN_38 = io_out_ready ? cmd_temp_pfch_tag : 7'h0; // @[CheckSplit.scala 186:51 CheckSplit.scala 143:33]
  wire [63:0] _GEN_43 = io_out_ready ? mini_addr : 64'h0; // @[CheckSplit.scala 186:51 CheckSplit.scala 143:33]
  wire [2:0] _GEN_44 = io_out_ready ? _GEN_32 : state; // @[CheckSplit.scala 186:51 CheckSplit.scala 138:28]
  wire  _T_11 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_55 = _T_10 ? state : 3'h0; // @[CheckSplit.scala 207:66 CheckSplit.scala 138:28 CheckSplit.scala 219:81]
  wire [2:0] _GEN_67 = io_out_ready ? _GEN_55 : state; // @[CheckSplit.scala 205:51 CheckSplit.scala 138:28]
  wire [63:0] _GEN_69 = _T_11 ? _GEN_34 : mini_addr; // @[Conditional.scala 39:67 CheckSplit.scala 133:32]
  wire [31:0] _GEN_70 = _T_11 ? _GEN_35 : mini_len; // @[Conditional.scala 39:67 CheckSplit.scala 134:31]
  wire  _GEN_71 = _T_11 & io_out_ready; // @[Conditional.scala 39:67 CheckSplit.scala 142:25]
  wire [31:0] _GEN_72 = _T_11 ? _GEN_37 : 32'h0; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [6:0] _GEN_73 = _T_11 ? _GEN_38 : 7'h0; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [63:0] _GEN_78 = _T_11 ? _GEN_43 : 64'h0; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [2:0] _GEN_79 = _T_11 ? _GEN_67 : state; // @[Conditional.scala 39:67 CheckSplit.scala 138:28]
  wire [63:0] _GEN_81 = _T_8 ? _GEN_34 : _GEN_69; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_82 = _T_8 ? _GEN_35 : _GEN_70; // @[Conditional.scala 39:67]
  wire  _GEN_83 = _T_8 ? io_out_ready : _GEN_71; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_84 = _T_8 ? _GEN_37 : _GEN_72; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_85 = _T_8 ? _GEN_38 : _GEN_73; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_90 = _T_8 ? _GEN_43 : _GEN_78; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_91 = _T_8 ? _GEN_44 : _GEN_79; // @[Conditional.scala 39:67]
  wire  _GEN_98 = _T_6 ? 1'h0 : _GEN_83; // @[Conditional.scala 39:67 CheckSplit.scala 142:25]
  wire [31:0] _GEN_99 = _T_6 ? 32'h0 : _GEN_84; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [6:0] _GEN_100 = _T_6 ? 7'h0 : _GEN_85; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [63:0] _GEN_105 = _T_6 ? 64'h0 : _GEN_90; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire  _GEN_112 = _T_2 ? 1'h0 : _GEN_98; // @[Conditional.scala 39:67 CheckSplit.scala 142:25]
  wire [31:0] _GEN_113 = _T_2 ? 32'h0 : _GEN_99; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [6:0] _GEN_114 = _T_2 ? 7'h0 : _GEN_100; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [63:0] _GEN_119 = _T_2 ? 64'h0 : _GEN_105; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [63:0] _GEN_129 = _T ? _GEN_9 : {{40'd0}, offset_addr}; // @[Conditional.scala 40:58 CheckSplit.scala 129:34]
  wire [63:0] _GEN_131 = _T ? _GEN_11 : {{40'd0}, new_length}; // @[Conditional.scala 40:58 CheckSplit.scala 130:33]
  assign io_in_ready = state == 3'h0; // @[CheckSplit.scala 140:35]
  assign io_out_valid = _T ? 1'h0 : _GEN_112; // @[Conditional.scala 40:58 CheckSplit.scala 142:25]
  assign io_out_bits_addr = _T ? 64'h0 : _GEN_119; // @[Conditional.scala 40:58 CheckSplit.scala 143:33]
  assign io_out_bits_pfch_tag = _T ? 7'h0 : _GEN_114; // @[Conditional.scala 40:58 CheckSplit.scala 143:33]
  assign io_out_bits_len = _T ? 32'h0 : _GEN_113; // @[Conditional.scala 40:58 CheckSplit.scala 143:33]
  always @(posedge clock) begin
    if (reset) begin // @[CheckSplit.scala 129:34]
      offset_addr <= 24'h0; // @[CheckSplit.scala 129:34]
    end else begin
      offset_addr <= _GEN_129[23:0];
    end
    if (reset) begin // @[CheckSplit.scala 130:33]
      new_length <= 24'h0; // @[CheckSplit.scala 130:33]
    end else begin
      new_length <= _GEN_131[23:0];
    end
    if (reset) begin // @[CheckSplit.scala 131:31]
      cmd_addr <= 64'h0; // @[CheckSplit.scala 131:31]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 150:43]
        cmd_addr <= io_in_bits_addr; // @[CheckSplit.scala 151:81]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 160:68]
        cmd_addr <= _cmd_addr_T_1; // @[CheckSplit.scala 163:81]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      cmd_addr <= _GEN_19;
    end
    if (reset) begin // @[CheckSplit.scala 132:30]
      cmd_len <= 32'h0; // @[CheckSplit.scala 132:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 150:43]
        cmd_len <= io_in_bits_len; // @[CheckSplit.scala 152:81]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 160:68]
        cmd_len <= _cmd_len_T_1; // @[CheckSplit.scala 164:81]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      cmd_len <= _GEN_20;
    end
    if (reset) begin // @[CheckSplit.scala 133:32]
      mini_addr <= 64'h0; // @[CheckSplit.scala 133:32]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        mini_addr <= cmd_addr;
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        mini_addr <= cmd_addr;
      end else begin
        mini_addr <= _GEN_81;
      end
    end
    if (reset) begin // @[CheckSplit.scala 134:31]
      mini_len <= 32'h0; // @[CheckSplit.scala 134:31]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 160:68]
          mini_len <= {{8'd0}, new_length}; // @[CheckSplit.scala 162:81]
        end else begin
          mini_len <= cmd_len; // @[CheckSplit.scala 168:81]
        end
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        mini_len <= _GEN_18;
      end else begin
        mini_len <= _GEN_82;
      end
    end
    if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 150:43]
        cmd_temp_pfch_tag <= io_in_bits_pfch_tag; // @[CheckSplit.scala 153:81]
      end
    end
    if (reset) begin // @[CheckSplit.scala 138:28]
      state <= 3'h0; // @[CheckSplit.scala 138:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 150:43]
        state <= 3'h1; // @[CheckSplit.scala 155:49]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 160:68]
        state <= 3'h3; // @[CheckSplit.scala 165:65]
      end else begin
        state <= 3'h4; // @[CheckSplit.scala 169:65]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      state <= _GEN_21;
    end else begin
      state <= _GEN_91;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_addr = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  new_length = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  cmd_addr = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  cmd_len = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  mini_addr = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  mini_len = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cmd_temp_pfch_tag = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CMDBoundaryCheck_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [31:0] io_in_bits_len,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [31:0] io_out_bits_len,
  output        io_out_bits_eop,
  output        io_out_bits_sop
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [23:0] offset_addr; // @[CheckSplit.scala 129:34]
  reg [23:0] new_length; // @[CheckSplit.scala 130:33]
  reg [63:0] cmd_addr; // @[CheckSplit.scala 131:31]
  reg [31:0] cmd_len; // @[CheckSplit.scala 132:30]
  reg [63:0] mini_addr; // @[CheckSplit.scala 133:32]
  reg [31:0] mini_len; // @[CheckSplit.scala 134:31]
  reg [2:0] state; // @[CheckSplit.scala 138:28]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _offset_addr_T = io_in_bits_addr & 64'h1fffff; // @[CheckSplit.scala 154:100]
  wire [63:0] _new_length_T_2 = 64'h200000 - _offset_addr_T; // @[CheckSplit.scala 156:96]
  wire [63:0] _GEN_14 = _T_1 ? _offset_addr_T : {{40'd0}, offset_addr}; // @[CheckSplit.scala 150:43 CheckSplit.scala 154:81 CheckSplit.scala 129:34]
  wire [63:0] _GEN_16 = _T_1 ? _new_length_T_2 : {{40'd0}, new_length}; // @[CheckSplit.scala 150:43 CheckSplit.scala 156:81 CheckSplit.scala 130:33]
  wire  _T_2 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_198 = {{8'd0}, offset_addr}; // @[CheckSplit.scala 160:43]
  wire [31:0] _T_4 = _GEN_198 + cmd_len; // @[CheckSplit.scala 160:43]
  wire [63:0] _GEN_199 = {{40'd0}, new_length}; // @[CheckSplit.scala 163:93]
  wire [63:0] _cmd_addr_T_1 = cmd_addr + _GEN_199; // @[CheckSplit.scala 163:93]
  wire [31:0] _GEN_200 = {{8'd0}, new_length}; // @[CheckSplit.scala 164:92]
  wire [31:0] _cmd_len_T_1 = cmd_len - _GEN_200; // @[CheckSplit.scala 164:92]
  wire  _T_6 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [63:0] _cmd_addr_T_3 = cmd_addr + 64'h200000; // @[CheckSplit.scala 176:93]
  wire [31:0] _cmd_len_T_3 = cmd_len - 32'h200000; // @[CheckSplit.scala 177:92]
  wire [31:0] _GEN_23 = cmd_len > 32'h200000 ? 32'h200000 : cmd_len; // @[CheckSplit.scala 173:52 CheckSplit.scala 175:81 CheckSplit.scala 181:81]
  wire [63:0] _GEN_24 = cmd_len > 32'h200000 ? _cmd_addr_T_3 : cmd_addr; // @[CheckSplit.scala 173:52 CheckSplit.scala 176:81 CheckSplit.scala 131:31]
  wire [31:0] _GEN_25 = cmd_len > 32'h200000 ? _cmd_len_T_3 : cmd_len; // @[CheckSplit.scala 173:52 CheckSplit.scala 177:81 CheckSplit.scala 132:30]
  wire [2:0] _GEN_26 = cmd_len > 32'h200000 ? 3'h3 : 3'h4; // @[CheckSplit.scala 173:52 CheckSplit.scala 178:65 CheckSplit.scala 182:65]
  wire  _T_8 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = mini_len > 32'h8000; // @[CheckSplit.scala 188:47]
  wire [63:0] _mini_addr_T_1 = mini_addr + 64'h8000; // @[CheckSplit.scala 189:94]
  wire [31:0] _mini_len_T_1 = mini_len - 32'h8000; // @[CheckSplit.scala 190:93]
  wire [63:0] _GEN_27 = mini_len > 32'h8000 ? _mini_addr_T_1 : mini_addr; // @[CheckSplit.scala 188:66 CheckSplit.scala 189:81 CheckSplit.scala 133:32]
  wire [31:0] _GEN_28 = mini_len > 32'h8000 ? _mini_len_T_1 : mini_len; // @[CheckSplit.scala 188:66 CheckSplit.scala 190:81 CheckSplit.scala 134:31]
  wire [31:0] _GEN_40 = mini_len > 32'h8000 ? 32'h8000 : mini_len; // @[CheckSplit.scala 188:66 CheckSplit.scala 193:73 CheckSplit.scala 198:73]
  wire [2:0] _GEN_42 = mini_len > 32'h8000 ? state : 3'h2; // @[CheckSplit.scala 188:66 CheckSplit.scala 138:28 CheckSplit.scala 200:81]
  wire [63:0] _GEN_44 = io_out_ready ? _GEN_27 : mini_addr; // @[CheckSplit.scala 186:51 CheckSplit.scala 133:32]
  wire [31:0] _GEN_45 = io_out_ready ? _GEN_28 : mini_len; // @[CheckSplit.scala 186:51 CheckSplit.scala 134:31]
  wire [31:0] _GEN_57 = io_out_ready ? _GEN_40 : 32'h0; // @[CheckSplit.scala 186:51 CheckSplit.scala 143:33]
  wire [63:0] _GEN_58 = io_out_ready ? mini_addr : 64'h0; // @[CheckSplit.scala 186:51 CheckSplit.scala 143:33]
  wire [2:0] _GEN_59 = io_out_ready ? _GEN_42 : state; // @[CheckSplit.scala 186:51 CheckSplit.scala 138:28]
  wire  _T_11 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_75 = _T_10 ? state : 3'h0; // @[CheckSplit.scala 207:66 CheckSplit.scala 138:28 CheckSplit.scala 219:81]
  wire [2:0] _GEN_92 = io_out_ready ? _GEN_75 : state; // @[CheckSplit.scala 205:51 CheckSplit.scala 138:28]
  wire [63:0] _GEN_94 = _T_11 ? _GEN_44 : mini_addr; // @[Conditional.scala 39:67 CheckSplit.scala 133:32]
  wire [31:0] _GEN_95 = _T_11 ? _GEN_45 : mini_len; // @[Conditional.scala 39:67 CheckSplit.scala 134:31]
  wire  _GEN_96 = _T_11 & io_out_ready; // @[Conditional.scala 39:67 CheckSplit.scala 142:25]
  wire [31:0] _GEN_107 = _T_11 ? _GEN_57 : 32'h0; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [63:0] _GEN_108 = _T_11 ? _GEN_58 : 64'h0; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [2:0] _GEN_109 = _T_11 ? _GEN_92 : state; // @[Conditional.scala 39:67 CheckSplit.scala 138:28]
  wire [63:0] _GEN_111 = _T_8 ? _GEN_44 : _GEN_94; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_112 = _T_8 ? _GEN_45 : _GEN_95; // @[Conditional.scala 39:67]
  wire  _GEN_113 = _T_8 ? io_out_ready : _GEN_96; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_124 = _T_8 ? _GEN_57 : _GEN_107; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_125 = _T_8 ? _GEN_58 : _GEN_108; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_126 = _T_8 ? _GEN_59 : _GEN_109; // @[Conditional.scala 39:67]
  wire  _GEN_133 = _T_6 ? 1'h0 : _GEN_113; // @[Conditional.scala 39:67 CheckSplit.scala 142:25]
  wire [31:0] _GEN_144 = _T_6 ? 32'h0 : _GEN_124; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [63:0] _GEN_145 = _T_6 ? 64'h0 : _GEN_125; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire  _GEN_152 = _T_2 ? 1'h0 : _GEN_133; // @[Conditional.scala 39:67 CheckSplit.scala 142:25]
  wire [31:0] _GEN_163 = _T_2 ? 32'h0 : _GEN_144; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [63:0] _GEN_164 = _T_2 ? 64'h0 : _GEN_145; // @[Conditional.scala 39:67 CheckSplit.scala 143:33]
  wire [63:0] _GEN_179 = _T ? _GEN_14 : {{40'd0}, offset_addr}; // @[Conditional.scala 40:58 CheckSplit.scala 129:34]
  wire [63:0] _GEN_181 = _T ? _GEN_16 : {{40'd0}, new_length}; // @[Conditional.scala 40:58 CheckSplit.scala 130:33]
  assign io_in_ready = state == 3'h0; // @[CheckSplit.scala 140:35]
  assign io_out_valid = _T ? 1'h0 : _GEN_152; // @[Conditional.scala 40:58 CheckSplit.scala 142:25]
  assign io_out_bits_addr = _T ? 64'h0 : _GEN_164; // @[Conditional.scala 40:58 CheckSplit.scala 143:33]
  assign io_out_bits_len = _T ? 32'h0 : _GEN_163; // @[Conditional.scala 40:58 CheckSplit.scala 143:33]
  assign io_out_bits_eop = _T ? 1'h0 : _GEN_152; // @[Conditional.scala 40:58 CheckSplit.scala 143:33]
  assign io_out_bits_sop = _T ? 1'h0 : _GEN_152; // @[Conditional.scala 40:58 CheckSplit.scala 143:33]
  always @(posedge clock) begin
    if (reset) begin // @[CheckSplit.scala 129:34]
      offset_addr <= 24'h0; // @[CheckSplit.scala 129:34]
    end else begin
      offset_addr <= _GEN_179[23:0];
    end
    if (reset) begin // @[CheckSplit.scala 130:33]
      new_length <= 24'h0; // @[CheckSplit.scala 130:33]
    end else begin
      new_length <= _GEN_181[23:0];
    end
    if (reset) begin // @[CheckSplit.scala 131:31]
      cmd_addr <= 64'h0; // @[CheckSplit.scala 131:31]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 150:43]
        cmd_addr <= io_in_bits_addr; // @[CheckSplit.scala 151:81]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 160:68]
        cmd_addr <= _cmd_addr_T_1; // @[CheckSplit.scala 163:81]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      cmd_addr <= _GEN_24;
    end
    if (reset) begin // @[CheckSplit.scala 132:30]
      cmd_len <= 32'h0; // @[CheckSplit.scala 132:30]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 150:43]
        cmd_len <= io_in_bits_len; // @[CheckSplit.scala 152:81]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 160:68]
        cmd_len <= _cmd_len_T_1; // @[CheckSplit.scala 164:81]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      cmd_len <= _GEN_25;
    end
    if (reset) begin // @[CheckSplit.scala 133:32]
      mini_addr <= 64'h0; // @[CheckSplit.scala 133:32]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        mini_addr <= cmd_addr;
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        mini_addr <= cmd_addr;
      end else begin
        mini_addr <= _GEN_111;
      end
    end
    if (reset) begin // @[CheckSplit.scala 134:31]
      mini_len <= 32'h0; // @[CheckSplit.scala 134:31]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[Conditional.scala 39:67]
        if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 160:68]
          mini_len <= {{8'd0}, new_length}; // @[CheckSplit.scala 162:81]
        end else begin
          mini_len <= cmd_len; // @[CheckSplit.scala 168:81]
        end
      end else if (_T_6) begin // @[Conditional.scala 39:67]
        mini_len <= _GEN_23;
      end else begin
        mini_len <= _GEN_112;
      end
    end
    if (reset) begin // @[CheckSplit.scala 138:28]
      state <= 3'h0; // @[CheckSplit.scala 138:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[CheckSplit.scala 150:43]
        state <= 3'h1; // @[CheckSplit.scala 155:49]
      end
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      if (_T_4 > 32'h200000) begin // @[CheckSplit.scala 160:68]
        state <= 3'h3; // @[CheckSplit.scala 165:65]
      end else begin
        state <= 3'h4; // @[CheckSplit.scala 169:65]
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      state <= _GEN_26;
    end else begin
      state <= _GEN_126;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  offset_addr = _RAND_0[23:0];
  _RAND_1 = {1{`RANDOM}};
  new_length = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  cmd_addr = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  cmd_len = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  mini_addr = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  mini_len = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XRam(
  input         clock,
  input         reset,
  input  [13:0] io_addr_a,
  input  [13:0] io_addr_b,
  input         io_wr_en_a,
  input  [63:0] io_data_in_a,
  output [63:0] io_data_out_a,
  output [63:0] io_data_out_b
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] ram_douta; // @[XRam.scala 136:33]
  wire [63:0] ram_doutb; // @[XRam.scala 136:33]
  wire [13:0] ram_addra; // @[XRam.scala 136:33]
  wire [13:0] ram_addrb; // @[XRam.scala 136:33]
  wire  ram_clka; // @[XRam.scala 136:33]
  wire  ram_clkb; // @[XRam.scala 136:33]
  wire [63:0] ram_dina; // @[XRam.scala 136:33]
  wire [63:0] ram_dinb; // @[XRam.scala 136:33]
  wire  ram_ena; // @[XRam.scala 136:33]
  wire  ram_enb; // @[XRam.scala 136:33]
  wire  ram_injectdbiterra; // @[XRam.scala 136:33]
  wire  ram_injectdbiterrb; // @[XRam.scala 136:33]
  wire  ram_injectsbiterra; // @[XRam.scala 136:33]
  wire  ram_injectsbiterrb; // @[XRam.scala 136:33]
  wire  ram_regcea; // @[XRam.scala 136:33]
  wire  ram_regceb; // @[XRam.scala 136:33]
  wire  ram_rsta; // @[XRam.scala 136:33]
  wire  ram_rstb; // @[XRam.scala 136:33]
  wire  ram_sleep; // @[XRam.scala 136:33]
  wire [7:0] ram_wea; // @[XRam.scala 136:33]
  wire [7:0] ram_web; // @[XRam.scala 136:33]
  wire [7:0] wr_en_a = io_wr_en_a ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  reg  usr_rst_delay_r; // @[Reg.scala 15:16]
  reg  usr_rst_delay_r_1; // @[Reg.scala 15:16]
  reg  usr_rst_delay_r_2; // @[Reg.scala 15:16]
  reg  usr_rst_delay; // @[Reg.scala 15:16]
  reg [13:0] reset_addr; // @[XRam.scala 141:54]
  wire [13:0] _reset_addr_T_1 = reset_addr + 14'h1; // @[XRam.scala 144:70]
  reg [13:0] r; // @[Reg.scala 15:16]
  reg [13:0] r_1; // @[Reg.scala 15:16]
  reg [13:0] REG; // @[XRam.scala 165:74]
  reg  REG_1; // @[XRam.scala 165:95]
  reg [63:0] io_data_out_b_REG; // @[XRam.scala 166:75]
  reg [13:0] r_2; // @[Reg.scala 15:16]
  reg [13:0] r_3; // @[Reg.scala 15:16]
  reg [13:0] r_4; // @[Reg.scala 15:16]
  reg [13:0] r_5; // @[Reg.scala 15:16]
  reg  r_6; // @[Reg.scala 15:16]
  reg  r_7; // @[Reg.scala 15:16]
  reg [63:0] io_data_out_b_r; // @[Reg.scala 15:16]
  reg [63:0] io_data_out_b_r_1; // @[Reg.scala 15:16]
  wire [63:0] _io_data_out_b_WIRE = ram_doutb; // @[XRam.scala 170:89 XRam.scala 170:89]
  wire [63:0] _GEN_15 = r_3 == r_5 & r_7 ? io_data_out_b_r_1 : _io_data_out_b_WIRE; // @[XRam.scala 167:130 XRam.scala 168:65 XRam.scala 170:65]
  xpm_memory_tdpram
    #(.USE_EMBEDDED_CONSTRAINT(0), .CLOCKING_MODE("common_clock"), .WRITE_DATA_WIDTH_B(64), .READ_LATENCY_B(2), .ADDR_WIDTH_A(14), .READ_DATA_WIDTH_A(64), .RST_MODE_B("SYNC"), .WAKEUP_TIME("disable_sleep"), .MEMORY_INIT_FILE("none"), .READ_LATENCY_A(2), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_A(64), .AUTO_SLEEP_TIME(0), .WRITE_MODE_A("no_change"), .MEMORY_PRIMITIVE("auto"), .USE_MEM_INIT(1), .MEMORY_INIT_PARAM(""), .SIM_ASSERT_CHK(0), .ECC_MODE("no_ecc"), .READ_RESET_VALUE_A("0"), .BYTE_WRITE_WIDTH_A(8), .MEMORY_OPTIMIZATION("true"), .MESSAGE_CONTROL(0), .WRITE_MODE_B("no_change"), .READ_DATA_WIDTH_B(64), .ADDR_WIDTH_B(14), .CASCADE_HEIGHT(0), .READ_RESET_VALUE_B("0"), .BYTE_WRITE_WIDTH_B(8), .MEMORY_SIZE(1048576))
    ram ( // @[XRam.scala 136:33]
    .douta(ram_douta),
    .doutb(ram_doutb),
    .addra(ram_addra),
    .addrb(ram_addrb),
    .clka(ram_clka),
    .clkb(ram_clkb),
    .dina(ram_dina),
    .dinb(ram_dinb),
    .ena(ram_ena),
    .enb(ram_enb),
    .injectdbiterra(ram_injectdbiterra),
    .injectdbiterrb(ram_injectdbiterrb),
    .injectsbiterra(ram_injectsbiterra),
    .injectsbiterrb(ram_injectsbiterrb),
    .regcea(ram_regcea),
    .regceb(ram_regceb),
    .rsta(ram_rsta),
    .rstb(ram_rstb),
    .sleep(ram_sleep),
    .wea(ram_wea),
    .web(ram_web)
  );
  assign io_data_out_a = ram_douta; // @[XRam.scala 175:73 XRam.scala 175:73]
  assign io_data_out_b = r_1 == REG & REG_1 ? io_data_out_b_REG : _GEN_15; // @[XRam.scala 165:108 XRam.scala 166:65]
  assign ram_addra = usr_rst_delay ? reset_addr : io_addr_a; // @[XRam.scala 178:55]
  assign ram_addrb = io_addr_b; // @[XRam.scala 179:49]
  assign ram_clka = clock; // @[XRam.scala 181:57]
  assign ram_clkb = clock; // @[XRam.scala 182:57]
  assign ram_dina = usr_rst_delay ? 64'h0 : io_data_in_a; // @[XRam.scala 184:63]
  assign ram_dinb = 64'h0; // @[XRam.scala 185:57]
  assign ram_ena = 1'h1; // @[XRam.scala 187:57]
  assign ram_enb = 1'h1; // @[XRam.scala 188:57]
  assign ram_injectdbiterra = 1'h0; // @[XRam.scala 190:41]
  assign ram_injectdbiterrb = 1'h0; // @[XRam.scala 191:41]
  assign ram_injectsbiterra = 1'h0; // @[XRam.scala 193:41]
  assign ram_injectsbiterrb = 1'h0; // @[XRam.scala 194:41]
  assign ram_regcea = 1'h1; // @[XRam.scala 196:49]
  assign ram_regceb = 1'h1; // @[XRam.scala 197:49]
  assign ram_rsta = 1'h0; // @[XRam.scala 199:57]
  assign ram_rstb = 1'h0; // @[XRam.scala 200:57]
  assign ram_sleep = 1'h0; // @[XRam.scala 202:49]
  assign ram_wea = usr_rst_delay ? 8'hff : wr_en_a; // @[XRam.scala 206:63]
  assign ram_web = 8'h0; // @[XRam.scala 208:57]
  always @(posedge clock) begin
    usr_rst_delay_r <= reset; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay_r_1 <= usr_rst_delay_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay_r_2 <= usr_rst_delay_r_1; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    usr_rst_delay <= usr_rst_delay_r_2; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    if (usr_rst_delay) begin // @[XRam.scala 143:45]
      reset_addr <= _reset_addr_T_1; // @[XRam.scala 144:57]
    end else begin
      reset_addr <= 14'h0; // @[XRam.scala 146:57]
    end
    r <= io_addr_b; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_1 <= r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    REG <= io_addr_a; // @[XRam.scala 165:74]
    REG_1 <= io_wr_en_a; // @[XRam.scala 165:95]
    io_data_out_b_REG <= io_data_in_a; // @[XRam.scala 166:75]
    r_2 <= io_addr_b; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_3 <= r_2; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_4 <= io_addr_a; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_5 <= r_4; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_6 <= io_wr_en_a; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    r_7 <= r_6; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    io_data_out_b_r <= io_data_in_a; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
    io_data_out_b_r_1 <= io_data_out_b_r; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  usr_rst_delay_r = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  usr_rst_delay_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  usr_rst_delay_r_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  usr_rst_delay = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  reset_addr = _RAND_4[13:0];
  _RAND_5 = {1{`RANDOM}};
  r = _RAND_5[13:0];
  _RAND_6 = {1{`RANDOM}};
  r_1 = _RAND_6[13:0];
  _RAND_7 = {1{`RANDOM}};
  REG = _RAND_7[13:0];
  _RAND_8 = {1{`RANDOM}};
  REG_1 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  io_data_out_b_REG = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  r_2 = _RAND_10[13:0];
  _RAND_11 = {1{`RANDOM}};
  r_3 = _RAND_11[13:0];
  _RAND_12 = {1{`RANDOM}};
  r_4 = _RAND_12[13:0];
  _RAND_13 = {1{`RANDOM}};
  r_5 = _RAND_13[13:0];
  _RAND_14 = {1{`RANDOM}};
  r_6 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  r_7 = _RAND_15[0:0];
  _RAND_16 = {2{`RANDOM}};
  io_data_out_b_r = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  io_data_out_b_r_1 = _RAND_17[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_addr,
  input  [31:0] io_enq_bits_len,
  input         io_enq_bits_eop,
  input         io_enq_bits_sop,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_addr,
  output [31:0] io_deq_bits_len,
  output        io_deq_bits_eop,
  output        io_deq_bits_sop,
  output        io_deq_bits_mrkr_req,
  output        io_deq_bits_sdi,
  output [10:0] io_deq_bits_qid,
  output        io_deq_bits_error,
  output [7:0]  io_deq_bits_func,
  output [15:0] io_deq_bits_cidx,
  output [2:0]  io_deq_bits_port_id,
  output        io_deq_bits_no_dma,
  output [3:0]  io_count
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_addr [0:9]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_len [0:9]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_eop [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_eop_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_eop_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_eop_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_eop_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_eop_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_eop_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_sop [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_sop_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_sop_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sop_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_sop_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sop_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_sop_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_mrkr_req [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_mrkr_req_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mrkr_req_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_mrkr_req_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mrkr_req_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_mrkr_req_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_mrkr_req_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_sdi [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_sdi_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_sdi_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sdi_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_sdi_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_sdi_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_sdi_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] ram_qid [0:9]; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_error [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_func [0:9]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_en; // @[Decoupled.scala 218:16]
  reg [15:0] ram_cidx [0:9]; // @[Decoupled.scala 218:16]
  wire [15:0] ram_cidx_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_cidx_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [15:0] ram_cidx_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_cidx_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_cidx_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_cidx_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_port_id [0:9]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_no_dma [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_no_dma_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_no_dma_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_no_dma_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_no_dma_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_no_dma_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_no_dma_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 4'h9; // @[Counter.scala 72:24]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire  wrap_1 = deq_ptr_value == 4'h9; // @[Counter.scala 72:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 257:32]
  wire [3:0] _io_count_T = maybe_full ? 4'ha : 4'h0; // @[Decoupled.scala 262:24]
  wire [3:0] _io_count_T_3 = 4'ha + ptr_diff; // @[Decoupled.scala 265:38]
  wire [3:0] _io_count_T_4 = deq_ptr_value > enq_ptr_value ? _io_count_T_3 : ptr_diff; // @[Decoupled.scala 264:24]
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_1[63:0] :
    ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_len_io_deq_bits_MPORT_data = ram_len_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_3[31:0] :
    ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_eop_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_eop_io_deq_bits_MPORT_data = ram_eop[ram_eop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_eop_io_deq_bits_MPORT_data = ram_eop_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_5[0:0] :
    ram_eop[ram_eop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_eop_MPORT_data = io_enq_bits_eop;
  assign ram_eop_MPORT_addr = enq_ptr_value;
  assign ram_eop_MPORT_mask = 1'h1;
  assign ram_eop_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sop_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_sop_io_deq_bits_MPORT_data = ram_sop[ram_sop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_sop_io_deq_bits_MPORT_data = ram_sop_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_7[0:0] :
    ram_sop[ram_sop_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_sop_MPORT_data = io_enq_bits_sop;
  assign ram_sop_MPORT_addr = enq_ptr_value;
  assign ram_sop_MPORT_mask = 1'h1;
  assign ram_sop_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mrkr_req_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mrkr_req_io_deq_bits_MPORT_data = ram_mrkr_req[ram_mrkr_req_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_mrkr_req_io_deq_bits_MPORT_data = ram_mrkr_req_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_9[0:0] :
    ram_mrkr_req[ram_mrkr_req_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_mrkr_req_MPORT_data = 1'h0;
  assign ram_mrkr_req_MPORT_addr = enq_ptr_value;
  assign ram_mrkr_req_MPORT_mask = 1'h1;
  assign ram_mrkr_req_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_sdi_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_sdi_io_deq_bits_MPORT_data = ram_sdi[ram_sdi_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_sdi_io_deq_bits_MPORT_data = ram_sdi_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_11[0:0] :
    ram_sdi[ram_sdi_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_sdi_MPORT_data = 1'h0;
  assign ram_sdi_MPORT_addr = enq_ptr_value;
  assign ram_sdi_MPORT_mask = 1'h1;
  assign ram_sdi_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qid_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_13[10:0] :
    ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_qid_MPORT_data = 11'h0;
  assign ram_qid_MPORT_addr = enq_ptr_value;
  assign ram_qid_MPORT_mask = 1'h1;
  assign ram_qid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_error_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_error_io_deq_bits_MPORT_data = ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_error_io_deq_bits_MPORT_data = ram_error_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_15[0:0] :
    ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_error_MPORT_data = 1'h0;
  assign ram_error_MPORT_addr = enq_ptr_value;
  assign ram_error_MPORT_mask = 1'h1;
  assign ram_error_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_func_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_func_io_deq_bits_MPORT_data = ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_func_io_deq_bits_MPORT_data = ram_func_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_17[7:0] :
    ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_func_MPORT_data = 8'h0;
  assign ram_func_MPORT_addr = enq_ptr_value;
  assign ram_func_MPORT_mask = 1'h1;
  assign ram_func_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_cidx_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_cidx_io_deq_bits_MPORT_data = ram_cidx[ram_cidx_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_cidx_io_deq_bits_MPORT_data = ram_cidx_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_19[15:0] :
    ram_cidx[ram_cidx_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_cidx_MPORT_data = 16'h0;
  assign ram_cidx_MPORT_addr = enq_ptr_value;
  assign ram_cidx_MPORT_mask = 1'h1;
  assign ram_cidx_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_port_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_21[2:0] :
    ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_port_id_MPORT_data = 3'h0;
  assign ram_port_id_MPORT_addr = enq_ptr_value;
  assign ram_port_id_MPORT_mask = 1'h1;
  assign ram_port_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_no_dma_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_no_dma_io_deq_bits_MPORT_data = ram_no_dma[ram_no_dma_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_no_dma_io_deq_bits_MPORT_data = ram_no_dma_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_23[0:0] :
    ram_no_dma[ram_no_dma_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_no_dma_MPORT_data = 1'h0;
  assign ram_no_dma_MPORT_addr = enq_ptr_value;
  assign ram_no_dma_MPORT_mask = 1'h1;
  assign ram_no_dma_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_eop = ram_eop_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_sop = ram_sop_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_mrkr_req = ram_mrkr_req_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_sdi = ram_sdi_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_qid = ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_error = ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_func = ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_cidx = ram_cidx_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_port_id = ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_no_dma = ram_no_dma_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_count = ptr_match ? _io_count_T : _io_count_T_4; // @[Decoupled.scala 261:20]
  always @(posedge clock) begin
    if(ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_eop_MPORT_en & ram_eop_MPORT_mask) begin
      ram_eop[ram_eop_MPORT_addr] <= ram_eop_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_sop_MPORT_en & ram_sop_MPORT_mask) begin
      ram_sop[ram_sop_MPORT_addr] <= ram_sop_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_mrkr_req_MPORT_en & ram_mrkr_req_MPORT_mask) begin
      ram_mrkr_req[ram_mrkr_req_MPORT_addr] <= ram_mrkr_req_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_sdi_MPORT_en & ram_sdi_MPORT_mask) begin
      ram_sdi[ram_sdi_MPORT_addr] <= ram_sdi_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_qid_MPORT_en & ram_qid_MPORT_mask) begin
      ram_qid[ram_qid_MPORT_addr] <= ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_error_MPORT_en & ram_error_MPORT_mask) begin
      ram_error[ram_error_MPORT_addr] <= ram_error_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_func_MPORT_en & ram_func_MPORT_mask) begin
      ram_func[ram_func_MPORT_addr] <= ram_func_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_cidx_MPORT_en & ram_cidx_MPORT_mask) begin
      ram_cidx[ram_cidx_MPORT_addr] <= ram_cidx_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_port_id_MPORT_en & ram_port_id_MPORT_mask) begin
      ram_port_id[ram_port_id_MPORT_addr] <= ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_no_dma_MPORT_en & ram_no_dma_MPORT_mask) begin
      ram_no_dma[ram_no_dma_MPORT_addr] <= ram_no_dma_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      if (wrap) begin // @[Counter.scala 86:20]
        enq_ptr_value <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      if (wrap_1) begin // @[Counter.scala 86:20]
        deq_ptr_value <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
  _RAND_17 = {1{`RANDOM}};
  _RAND_19 = {1{`RANDOM}};
  _RAND_21 = {1{`RANDOM}};
  _RAND_23 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_len[initvar] = _RAND_2[31:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_eop[initvar] = _RAND_4[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_sop[initvar] = _RAND_6[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_mrkr_req[initvar] = _RAND_8[0:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_sdi[initvar] = _RAND_10[0:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_qid[initvar] = _RAND_12[10:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_error[initvar] = _RAND_14[0:0];
  _RAND_16 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_func[initvar] = _RAND_16[7:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_cidx[initvar] = _RAND_18[15:0];
  _RAND_20 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_port_id[initvar] = _RAND_20[2:0];
  _RAND_22 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_no_dma[initvar] = _RAND_22[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  enq_ptr_value = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  deq_ptr_value = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  maybe_full = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_1(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_addr,
  input  [6:0]  io_enq_bits_pfch_tag,
  input  [31:0] io_enq_bits_len,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_addr,
  output [10:0] io_deq_bits_qid,
  output        io_deq_bits_error,
  output [7:0]  io_deq_bits_func,
  output [2:0]  io_deq_bits_port_id,
  output [6:0]  io_deq_bits_pfch_tag,
  output [31:0] io_deq_bits_len,
  output [3:0]  io_count
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_addr [0:9]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] ram_qid [0:9]; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_error [0:9]; // @[Decoupled.scala 218:16]
  wire  ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_func [0:9]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_port_id [0:9]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_pfch_tag [0:9]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_pfch_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_pfch_tag_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_pfch_tag_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_pfch_tag_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_pfch_tag_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_pfch_tag_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_len [0:9]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire  wrap = enq_ptr_value == 4'h9; // @[Counter.scala 72:24]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire  wrap_1 = deq_ptr_value == 4'h9; // @[Counter.scala 72:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] ptr_diff = enq_ptr_value - deq_ptr_value; // @[Decoupled.scala 257:32]
  wire [3:0] _io_count_T = maybe_full ? 4'ha : 4'h0; // @[Decoupled.scala 262:24]
  wire [3:0] _io_count_T_3 = 4'ha + ptr_diff; // @[Decoupled.scala 265:38]
  wire [3:0] _io_count_T_4 = deq_ptr_value > enq_ptr_value ? _io_count_T_3 : ptr_diff; // @[Decoupled.scala 264:24]
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_1[63:0] :
    ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qid_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_3[10:0] :
    ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_qid_MPORT_data = 11'h0;
  assign ram_qid_MPORT_addr = enq_ptr_value;
  assign ram_qid_MPORT_mask = 1'h1;
  assign ram_qid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_error_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_error_io_deq_bits_MPORT_data = ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_error_io_deq_bits_MPORT_data = ram_error_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_5[0:0] :
    ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_error_MPORT_data = 1'h0;
  assign ram_error_MPORT_addr = enq_ptr_value;
  assign ram_error_MPORT_mask = 1'h1;
  assign ram_error_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_func_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_func_io_deq_bits_MPORT_data = ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_func_io_deq_bits_MPORT_data = ram_func_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_7[7:0] :
    ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_func_MPORT_data = 8'h0;
  assign ram_func_MPORT_addr = enq_ptr_value;
  assign ram_func_MPORT_mask = 1'h1;
  assign ram_func_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_port_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_9[2:0] :
    ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_port_id_MPORT_data = 3'h0;
  assign ram_port_id_MPORT_addr = enq_ptr_value;
  assign ram_port_id_MPORT_mask = 1'h1;
  assign ram_port_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pfch_tag_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_pfch_tag_io_deq_bits_MPORT_data = ram_pfch_tag[ram_pfch_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_pfch_tag_io_deq_bits_MPORT_data = ram_pfch_tag_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_11[6:0] :
    ram_pfch_tag[ram_pfch_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_pfch_tag_MPORT_data = io_enq_bits_pfch_tag;
  assign ram_pfch_tag_MPORT_addr = enq_ptr_value;
  assign ram_pfch_tag_MPORT_mask = 1'h1;
  assign ram_pfch_tag_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `else
  assign ram_len_io_deq_bits_MPORT_data = ram_len_io_deq_bits_MPORT_addr >= 4'ha ? _RAND_13[31:0] :
    ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_qid = ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_error = ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_func = ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_port_id = ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_pfch_tag = ram_pfch_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_count = ptr_match ? _io_count_T : _io_count_T_4; // @[Decoupled.scala 261:20]
  always @(posedge clock) begin
    if(ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_qid_MPORT_en & ram_qid_MPORT_mask) begin
      ram_qid[ram_qid_MPORT_addr] <= ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_error_MPORT_en & ram_error_MPORT_mask) begin
      ram_error[ram_error_MPORT_addr] <= ram_error_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_func_MPORT_en & ram_func_MPORT_mask) begin
      ram_func[ram_func_MPORT_addr] <= ram_func_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_port_id_MPORT_en & ram_port_id_MPORT_mask) begin
      ram_port_id[ram_port_id_MPORT_addr] <= ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_pfch_tag_MPORT_en & ram_pfch_tag_MPORT_mask) begin
      ram_pfch_tag[ram_pfch_tag_MPORT_addr] <= ram_pfch_tag_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      if (wrap) begin // @[Counter.scala 86:20]
        enq_ptr_value <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      if (wrap_1) begin // @[Counter.scala 86:20]
        deq_ptr_value <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[63:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_qid[initvar] = _RAND_2[10:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_error[initvar] = _RAND_4[0:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_func[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_port_id[initvar] = _RAND_8[2:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_pfch_tag[initvar] = _RAND_10[6:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 10; initvar = initvar+1)
    ram_len[initvar] = _RAND_12[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  enq_ptr_value = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  deq_ptr_value = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  maybe_full = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TLB(
  input         clock,
  input         reset,
  output        io_wr_tlb_ready,
  input         io_wr_tlb_valid,
  input  [31:0] io_wr_tlb_bits_vaddr_high,
  input  [31:0] io_wr_tlb_bits_vaddr_low,
  input  [31:0] io_wr_tlb_bits_paddr_high,
  input  [31:0] io_wr_tlb_bits_paddr_low,
  input         io_wr_tlb_bits_is_base,
  output        io_h2c_in_ready,
  input         io_h2c_in_valid,
  input  [63:0] io_h2c_in_bits_addr,
  input  [31:0] io_h2c_in_bits_len,
  input         io_h2c_in_bits_eop,
  input         io_h2c_in_bits_sop,
  output        io_c2h_in_ready,
  input         io_c2h_in_valid,
  input  [63:0] io_c2h_in_bits_addr,
  input  [6:0]  io_c2h_in_bits_pfch_tag,
  input  [31:0] io_c2h_in_bits_len,
  input         io_h2c_out_ready,
  output        io_h2c_out_valid,
  output [63:0] io_h2c_out_bits_addr,
  output [31:0] io_h2c_out_bits_len,
  output        io_h2c_out_bits_eop,
  output        io_h2c_out_bits_sop,
  output        io_h2c_out_bits_mrkr_req,
  output        io_h2c_out_bits_sdi,
  output [10:0] io_h2c_out_bits_qid,
  output        io_h2c_out_bits_error,
  output [7:0]  io_h2c_out_bits_func,
  output [15:0] io_h2c_out_bits_cidx,
  output [2:0]  io_h2c_out_bits_port_id,
  output        io_h2c_out_bits_no_dma,
  input         io_c2h_out_ready,
  output        io_c2h_out_valid,
  output [63:0] io_c2h_out_bits_addr,
  output [10:0] io_c2h_out_bits_qid,
  output        io_c2h_out_bits_error,
  output [7:0]  io_c2h_out_bits_func,
  output [2:0]  io_c2h_out_bits_port_id,
  output [6:0]  io_c2h_out_bits_pfch_tag,
  output [31:0] io_c2h_out_bits_len,
  output [31:0] io_tlb_miss_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  tlb_table_clock; // @[XRam.scala 102:23]
  wire  tlb_table_reset; // @[XRam.scala 102:23]
  wire [13:0] tlb_table_io_addr_a; // @[XRam.scala 102:23]
  wire [13:0] tlb_table_io_addr_b; // @[XRam.scala 102:23]
  wire  tlb_table_io_wr_en_a; // @[XRam.scala 102:23]
  wire [63:0] tlb_table_io_data_in_a; // @[XRam.scala 102:23]
  wire [63:0] tlb_table_io_data_out_a; // @[XRam.scala 102:23]
  wire [63:0] tlb_table_io_data_out_b; // @[XRam.scala 102:23]
  wire  q_h2c_clock; // @[TLB.scala 71:57]
  wire  q_h2c_reset; // @[TLB.scala 71:57]
  wire  q_h2c_io_enq_ready; // @[TLB.scala 71:57]
  wire  q_h2c_io_enq_valid; // @[TLB.scala 71:57]
  wire [63:0] q_h2c_io_enq_bits_addr; // @[TLB.scala 71:57]
  wire [31:0] q_h2c_io_enq_bits_len; // @[TLB.scala 71:57]
  wire  q_h2c_io_enq_bits_eop; // @[TLB.scala 71:57]
  wire  q_h2c_io_enq_bits_sop; // @[TLB.scala 71:57]
  wire  q_h2c_io_deq_ready; // @[TLB.scala 71:57]
  wire  q_h2c_io_deq_valid; // @[TLB.scala 71:57]
  wire [63:0] q_h2c_io_deq_bits_addr; // @[TLB.scala 71:57]
  wire [31:0] q_h2c_io_deq_bits_len; // @[TLB.scala 71:57]
  wire  q_h2c_io_deq_bits_eop; // @[TLB.scala 71:57]
  wire  q_h2c_io_deq_bits_sop; // @[TLB.scala 71:57]
  wire  q_h2c_io_deq_bits_mrkr_req; // @[TLB.scala 71:57]
  wire  q_h2c_io_deq_bits_sdi; // @[TLB.scala 71:57]
  wire [10:0] q_h2c_io_deq_bits_qid; // @[TLB.scala 71:57]
  wire  q_h2c_io_deq_bits_error; // @[TLB.scala 71:57]
  wire [7:0] q_h2c_io_deq_bits_func; // @[TLB.scala 71:57]
  wire [15:0] q_h2c_io_deq_bits_cidx; // @[TLB.scala 71:57]
  wire [2:0] q_h2c_io_deq_bits_port_id; // @[TLB.scala 71:57]
  wire  q_h2c_io_deq_bits_no_dma; // @[TLB.scala 71:57]
  wire [3:0] q_h2c_io_count; // @[TLB.scala 71:57]
  wire  q_c2h_clock; // @[TLB.scala 72:57]
  wire  q_c2h_reset; // @[TLB.scala 72:57]
  wire  q_c2h_io_enq_ready; // @[TLB.scala 72:57]
  wire  q_c2h_io_enq_valid; // @[TLB.scala 72:57]
  wire [63:0] q_c2h_io_enq_bits_addr; // @[TLB.scala 72:57]
  wire [6:0] q_c2h_io_enq_bits_pfch_tag; // @[TLB.scala 72:57]
  wire [31:0] q_c2h_io_enq_bits_len; // @[TLB.scala 72:57]
  wire  q_c2h_io_deq_ready; // @[TLB.scala 72:57]
  wire  q_c2h_io_deq_valid; // @[TLB.scala 72:57]
  wire [63:0] q_c2h_io_deq_bits_addr; // @[TLB.scala 72:57]
  wire [10:0] q_c2h_io_deq_bits_qid; // @[TLB.scala 72:57]
  wire  q_c2h_io_deq_bits_error; // @[TLB.scala 72:57]
  wire [7:0] q_c2h_io_deq_bits_func; // @[TLB.scala 72:57]
  wire [2:0] q_c2h_io_deq_bits_port_id; // @[TLB.scala 72:57]
  wire [6:0] q_c2h_io_deq_bits_pfch_tag; // @[TLB.scala 72:57]
  wire [31:0] q_c2h_io_deq_bits_len; // @[TLB.scala 72:57]
  wire [3:0] q_c2h_io_count; // @[TLB.scala 72:57]
  reg [42:0] base_page; // @[TLB.scala 33:50]
  reg [31:0] tlb_miss_count; // @[TLB.scala 34:50]
  reg [14:0] wrtlb_index; // @[TLB.scala 36:50]
  wire [42:0] h2c_page = io_h2c_in_bits_addr[63:21]; // @[TLB.scala 37:62]
  wire [42:0] h2c_index = h2c_page - base_page; // @[TLB.scala 38:52]
  wire [42:0] _GEN_12 = {{28'd0}, wrtlb_index}; // @[TLB.scala 39:90]
  wire [42:0] _h2c_outrange_T_2 = base_page + _GEN_12; // @[TLB.scala 39:90]
  wire  h2c_outrange = h2c_page < base_page | h2c_page >= _h2c_outrange_T_2; // @[TLB.scala 39:66]
  wire [42:0] c2h_page = io_c2h_in_bits_addr[63:21]; // @[TLB.scala 40:62]
  wire [42:0] c2h_index = c2h_page - base_page; // @[TLB.scala 41:52]
  wire  c2h_outrange = c2h_page < base_page | c2h_page >= _h2c_outrange_T_2; // @[TLB.scala 42:66]
  wire  _tlb_table_io_wr_en_a_T = io_wr_tlb_ready & io_wr_tlb_valid; // @[Decoupled.scala 40:37]
  wire [14:0] _wrtlb_index_T_1 = wrtlb_index + 15'h1; // @[TLB.scala 53:72]
  wire [63:0] _base_page_T = {io_wr_tlb_bits_vaddr_high,io_wr_tlb_bits_vaddr_low}; // @[Cat.scala 30:58]
  wire [14:0] _GEN_1 = io_wr_tlb_bits_is_base ? 15'h0 : wrtlb_index; // @[TLB.scala 54:51 TLB.scala 56:49 TLB.scala 52:49]
  wire [42:0] _GEN_4 = _tlb_table_io_wr_en_a_T ? {{28'd0}, _GEN_1} : h2c_index; // @[TLB.scala 51:31 TLB.scala 61:41]
  reg [31:0] h2c_bits_delay_REG_len; // @[TLB.scala 67:59]
  reg  h2c_bits_delay_REG_eop; // @[TLB.scala 67:59]
  reg  h2c_bits_delay_REG_sop; // @[TLB.scala 67:59]
  reg [31:0] h2c_bits_delay_REG_1_len; // @[TLB.scala 67:51]
  reg  h2c_bits_delay_REG_1_eop; // @[TLB.scala 67:51]
  reg  h2c_bits_delay_REG_1_sop; // @[TLB.scala 67:51]
  reg [6:0] c2h_bits_delay_REG_pfch_tag; // @[TLB.scala 68:59]
  reg [31:0] c2h_bits_delay_REG_len; // @[TLB.scala 68:59]
  reg [6:0] c2h_bits_delay_REG_1_pfch_tag; // @[TLB.scala 68:51]
  reg [31:0] c2h_bits_delay_REG_1_len; // @[TLB.scala 68:51]
  reg [20:0] h2c_bits_delay_addr_REG; // @[TLB.scala 69:77]
  reg [20:0] h2c_bits_delay_addr_REG_1; // @[TLB.scala 69:69]
  wire [63:0] _GEN_14 = {{43'd0}, h2c_bits_delay_addr_REG_1}; // @[TLB.scala 69:60]
  reg [20:0] c2h_bits_delay_addr_REG; // @[TLB.scala 70:77]
  reg [20:0] c2h_bits_delay_addr_REG_1; // @[TLB.scala 70:69]
  wire [63:0] _GEN_15 = {{43'd0}, c2h_bits_delay_addr_REG_1}; // @[TLB.scala 70:60]
  reg  REG; // @[TLB.scala 77:29]
  reg  REG_1; // @[TLB.scala 77:21]
  reg  REG_2; // @[TLB.scala 77:66]
  reg  REG_3; // @[TLB.scala 77:58]
  reg  REG_4; // @[TLB.scala 77:104]
  reg  REG_5; // @[TLB.scala 77:96]
  reg  REG_6; // @[TLB.scala 83:29]
  reg  REG_7; // @[TLB.scala 83:21]
  reg  REG_8; // @[TLB.scala 83:66]
  reg  REG_9; // @[TLB.scala 83:58]
  reg  REG_10; // @[TLB.scala 83:104]
  reg  REG_11; // @[TLB.scala 83:96]
  wire  h2c_miss = h2c_outrange & io_h2c_in_valid & io_h2c_in_ready; // @[TLB.scala 89:58]
  wire  c2h_miss = c2h_outrange & io_c2h_in_valid & io_c2h_in_ready; // @[TLB.scala 90:58]
  wire [31:0] _tlb_miss_count_T_1 = tlb_miss_count + 32'h1; // @[TLB.scala 92:50]
  wire [31:0] _tlb_miss_count_T_3 = tlb_miss_count + 32'h2; // @[TLB.scala 94:58]
  XRam tlb_table ( // @[XRam.scala 102:23]
    .clock(tlb_table_clock),
    .reset(tlb_table_reset),
    .io_addr_a(tlb_table_io_addr_a),
    .io_addr_b(tlb_table_io_addr_b),
    .io_wr_en_a(tlb_table_io_wr_en_a),
    .io_data_in_a(tlb_table_io_data_in_a),
    .io_data_out_a(tlb_table_io_data_out_a),
    .io_data_out_b(tlb_table_io_data_out_b)
  );
  Queue q_h2c ( // @[TLB.scala 71:57]
    .clock(q_h2c_clock),
    .reset(q_h2c_reset),
    .io_enq_ready(q_h2c_io_enq_ready),
    .io_enq_valid(q_h2c_io_enq_valid),
    .io_enq_bits_addr(q_h2c_io_enq_bits_addr),
    .io_enq_bits_len(q_h2c_io_enq_bits_len),
    .io_enq_bits_eop(q_h2c_io_enq_bits_eop),
    .io_enq_bits_sop(q_h2c_io_enq_bits_sop),
    .io_deq_ready(q_h2c_io_deq_ready),
    .io_deq_valid(q_h2c_io_deq_valid),
    .io_deq_bits_addr(q_h2c_io_deq_bits_addr),
    .io_deq_bits_len(q_h2c_io_deq_bits_len),
    .io_deq_bits_eop(q_h2c_io_deq_bits_eop),
    .io_deq_bits_sop(q_h2c_io_deq_bits_sop),
    .io_deq_bits_mrkr_req(q_h2c_io_deq_bits_mrkr_req),
    .io_deq_bits_sdi(q_h2c_io_deq_bits_sdi),
    .io_deq_bits_qid(q_h2c_io_deq_bits_qid),
    .io_deq_bits_error(q_h2c_io_deq_bits_error),
    .io_deq_bits_func(q_h2c_io_deq_bits_func),
    .io_deq_bits_cidx(q_h2c_io_deq_bits_cidx),
    .io_deq_bits_port_id(q_h2c_io_deq_bits_port_id),
    .io_deq_bits_no_dma(q_h2c_io_deq_bits_no_dma),
    .io_count(q_h2c_io_count)
  );
  Queue_1 q_c2h ( // @[TLB.scala 72:57]
    .clock(q_c2h_clock),
    .reset(q_c2h_reset),
    .io_enq_ready(q_c2h_io_enq_ready),
    .io_enq_valid(q_c2h_io_enq_valid),
    .io_enq_bits_addr(q_c2h_io_enq_bits_addr),
    .io_enq_bits_pfch_tag(q_c2h_io_enq_bits_pfch_tag),
    .io_enq_bits_len(q_c2h_io_enq_bits_len),
    .io_deq_ready(q_c2h_io_deq_ready),
    .io_deq_valid(q_c2h_io_deq_valid),
    .io_deq_bits_addr(q_c2h_io_deq_bits_addr),
    .io_deq_bits_qid(q_c2h_io_deq_bits_qid),
    .io_deq_bits_error(q_c2h_io_deq_bits_error),
    .io_deq_bits_func(q_c2h_io_deq_bits_func),
    .io_deq_bits_port_id(q_c2h_io_deq_bits_port_id),
    .io_deq_bits_pfch_tag(q_c2h_io_deq_bits_pfch_tag),
    .io_deq_bits_len(q_c2h_io_deq_bits_len),
    .io_count(q_c2h_io_count)
  );
  assign io_wr_tlb_ready = 1'h1; // @[TLB.scala 47:41]
  assign io_h2c_in_ready = q_h2c_io_count < 4'h8; // @[TLB.scala 74:59]
  assign io_c2h_in_ready = q_c2h_io_count < 4'h8; // @[TLB.scala 75:59]
  assign io_h2c_out_valid = q_h2c_io_deq_valid; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_addr = q_h2c_io_deq_bits_addr; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_len = q_h2c_io_deq_bits_len; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_eop = q_h2c_io_deq_bits_eop; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_sop = q_h2c_io_deq_bits_sop; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_mrkr_req = q_h2c_io_deq_bits_mrkr_req; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_sdi = q_h2c_io_deq_bits_sdi; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_qid = q_h2c_io_deq_bits_qid; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_error = q_h2c_io_deq_bits_error; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_func = q_h2c_io_deq_bits_func; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_cidx = q_h2c_io_deq_bits_cidx; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_port_id = q_h2c_io_deq_bits_port_id; // @[TLB.scala 99:41]
  assign io_h2c_out_bits_no_dma = q_h2c_io_deq_bits_no_dma; // @[TLB.scala 99:41]
  assign io_c2h_out_valid = q_c2h_io_deq_valid; // @[TLB.scala 102:41]
  assign io_c2h_out_bits_addr = q_c2h_io_deq_bits_addr; // @[TLB.scala 102:41]
  assign io_c2h_out_bits_qid = q_c2h_io_deq_bits_qid; // @[TLB.scala 102:41]
  assign io_c2h_out_bits_error = q_c2h_io_deq_bits_error; // @[TLB.scala 102:41]
  assign io_c2h_out_bits_func = q_c2h_io_deq_bits_func; // @[TLB.scala 102:41]
  assign io_c2h_out_bits_port_id = q_c2h_io_deq_bits_port_id; // @[TLB.scala 102:41]
  assign io_c2h_out_bits_pfch_tag = q_c2h_io_deq_bits_pfch_tag; // @[TLB.scala 102:41]
  assign io_c2h_out_bits_len = q_c2h_io_deq_bits_len; // @[TLB.scala 102:41]
  assign io_tlb_miss_count = tlb_miss_count; // @[TLB.scala 104:33]
  assign tlb_table_clock = clock;
  assign tlb_table_reset = reset;
  assign tlb_table_io_addr_a = _GEN_4[13:0];
  assign tlb_table_io_addr_b = c2h_index[13:0]; // @[TLB.scala 63:41]
  assign tlb_table_io_wr_en_a = io_wr_tlb_ready & io_wr_tlb_valid; // @[Decoupled.scala 40:37]
  assign tlb_table_io_data_in_a = {io_wr_tlb_bits_paddr_high,io_wr_tlb_bits_paddr_low}; // @[Cat.scala 30:58]
  assign q_h2c_clock = clock;
  assign q_h2c_reset = reset;
  assign q_h2c_io_enq_valid = REG_1 & REG_3 & ~REG_5; // @[TLB.scala 77:85]
  assign q_h2c_io_enq_bits_addr = tlb_table_io_data_out_a + _GEN_14; // @[TLB.scala 69:60]
  assign q_h2c_io_enq_bits_len = h2c_bits_delay_REG_1_len; // @[TLB.scala 65:47 TLB.scala 67:41]
  assign q_h2c_io_enq_bits_eop = h2c_bits_delay_REG_1_eop; // @[TLB.scala 65:47 TLB.scala 67:41]
  assign q_h2c_io_enq_bits_sop = h2c_bits_delay_REG_1_sop; // @[TLB.scala 65:47 TLB.scala 67:41]
  assign q_h2c_io_deq_ready = io_h2c_out_ready; // @[TLB.scala 99:41]
  assign q_c2h_clock = clock;
  assign q_c2h_reset = reset;
  assign q_c2h_io_enq_valid = REG_7 & REG_9 & ~REG_11; // @[TLB.scala 83:85]
  assign q_c2h_io_enq_bits_addr = tlb_table_io_data_out_b + _GEN_15; // @[TLB.scala 70:60]
  assign q_c2h_io_enq_bits_pfch_tag = c2h_bits_delay_REG_1_pfch_tag; // @[TLB.scala 66:47 TLB.scala 68:41]
  assign q_c2h_io_enq_bits_len = c2h_bits_delay_REG_1_len; // @[TLB.scala 66:47 TLB.scala 68:41]
  assign q_c2h_io_deq_ready = io_c2h_out_ready; // @[TLB.scala 102:41]
  always @(posedge clock) begin
    if (reset) begin // @[TLB.scala 33:50]
      base_page <= 43'h0; // @[TLB.scala 33:50]
    end else if (_tlb_table_io_wr_en_a_T) begin // @[TLB.scala 51:31]
      if (io_wr_tlb_bits_is_base) begin // @[TLB.scala 54:51]
        base_page <= _base_page_T[63:21]; // @[TLB.scala 55:57]
      end
    end
    if (reset) begin // @[TLB.scala 34:50]
      tlb_miss_count <= 32'h0; // @[TLB.scala 34:50]
    end else if (h2c_miss | c2h_miss) begin // @[TLB.scala 91:34]
      if (h2c_miss & c2h_miss) begin // @[TLB.scala 93:42]
        tlb_miss_count <= _tlb_miss_count_T_3; // @[TLB.scala 94:41]
      end else begin
        tlb_miss_count <= _tlb_miss_count_T_1; // @[TLB.scala 92:33]
      end
    end else if (_tlb_table_io_wr_en_a_T) begin // @[TLB.scala 51:31]
      if (io_wr_tlb_bits_is_base) begin // @[TLB.scala 54:51]
        tlb_miss_count <= 32'h0; // @[TLB.scala 58:49]
      end
    end
    if (reset) begin // @[TLB.scala 36:50]
      wrtlb_index <= 15'h0; // @[TLB.scala 36:50]
    end else if (_tlb_table_io_wr_en_a_T) begin // @[TLB.scala 51:31]
      if (io_wr_tlb_bits_is_base) begin // @[TLB.scala 54:51]
        wrtlb_index <= 15'h1; // @[TLB.scala 57:57]
      end else begin
        wrtlb_index <= _wrtlb_index_T_1; // @[TLB.scala 53:57]
      end
    end
    h2c_bits_delay_REG_len <= io_h2c_in_bits_len; // @[TLB.scala 67:59]
    h2c_bits_delay_REG_eop <= io_h2c_in_bits_eop; // @[TLB.scala 67:59]
    h2c_bits_delay_REG_sop <= io_h2c_in_bits_sop; // @[TLB.scala 67:59]
    h2c_bits_delay_REG_1_len <= h2c_bits_delay_REG_len; // @[TLB.scala 67:51]
    h2c_bits_delay_REG_1_eop <= h2c_bits_delay_REG_eop; // @[TLB.scala 67:51]
    h2c_bits_delay_REG_1_sop <= h2c_bits_delay_REG_sop; // @[TLB.scala 67:51]
    c2h_bits_delay_REG_pfch_tag <= io_c2h_in_bits_pfch_tag; // @[TLB.scala 68:59]
    c2h_bits_delay_REG_len <= io_c2h_in_bits_len; // @[TLB.scala 68:59]
    c2h_bits_delay_REG_1_pfch_tag <= c2h_bits_delay_REG_pfch_tag; // @[TLB.scala 68:51]
    c2h_bits_delay_REG_1_len <= c2h_bits_delay_REG_len; // @[TLB.scala 68:51]
    h2c_bits_delay_addr_REG <= io_h2c_in_bits_addr[20:0]; // @[TLB.scala 69:97]
    h2c_bits_delay_addr_REG_1 <= h2c_bits_delay_addr_REG; // @[TLB.scala 69:69]
    c2h_bits_delay_addr_REG <= io_c2h_in_bits_addr[20:0]; // @[TLB.scala 70:97]
    c2h_bits_delay_addr_REG_1 <= c2h_bits_delay_addr_REG; // @[TLB.scala 70:69]
    REG <= io_h2c_in_valid; // @[TLB.scala 77:29]
    REG_1 <= REG; // @[TLB.scala 77:21]
    REG_2 <= io_h2c_in_ready; // @[TLB.scala 77:66]
    REG_3 <= REG_2; // @[TLB.scala 77:58]
    REG_4 <= h2c_page < base_page | h2c_page >= _h2c_outrange_T_2; // @[TLB.scala 39:66]
    REG_5 <= REG_4; // @[TLB.scala 77:96]
    REG_6 <= io_c2h_in_valid; // @[TLB.scala 83:29]
    REG_7 <= REG_6; // @[TLB.scala 83:21]
    REG_8 <= io_c2h_in_ready; // @[TLB.scala 83:66]
    REG_9 <= REG_8; // @[TLB.scala 83:58]
    REG_10 <= c2h_page < base_page | c2h_page >= _h2c_outrange_T_2; // @[TLB.scala 42:66]
    REG_11 <= REG_10; // @[TLB.scala 83:96]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  base_page = _RAND_0[42:0];
  _RAND_1 = {1{`RANDOM}};
  tlb_miss_count = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  wrtlb_index = _RAND_2[14:0];
  _RAND_3 = {1{`RANDOM}};
  h2c_bits_delay_REG_len = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  h2c_bits_delay_REG_eop = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  h2c_bits_delay_REG_sop = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_len = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_eop = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  h2c_bits_delay_REG_1_sop = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  c2h_bits_delay_REG_pfch_tag = _RAND_9[6:0];
  _RAND_10 = {1{`RANDOM}};
  c2h_bits_delay_REG_len = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2h_bits_delay_REG_1_pfch_tag = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  c2h_bits_delay_REG_1_len = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  h2c_bits_delay_addr_REG = _RAND_13[20:0];
  _RAND_14 = {1{`RANDOM}};
  h2c_bits_delay_addr_REG_1 = _RAND_14[20:0];
  _RAND_15 = {1{`RANDOM}};
  c2h_bits_delay_addr_REG = _RAND_15[20:0];
  _RAND_16 = {1{`RANDOM}};
  c2h_bits_delay_addr_REG_1 = _RAND_16[20:0];
  _RAND_17 = {1{`RANDOM}};
  REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  REG_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  REG_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  REG_3 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  REG_4 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  REG_5 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  REG_6 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  REG_7 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  REG_8 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  REG_9 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  REG_10 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  REG_11 = _RAND_28[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SV_STREAM_FIFO_4(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [135:0] io_in_data,
  input          io_in_valid,
  output [135:0] io_out_data,
  output         io_out_valid
);
  wire [135:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [16:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [4:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [4:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [135:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [16:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [16:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(5), .CLOCKING_MODE("independent_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(16), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(5), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(136), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = 1'h1; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 17'h1ffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 17'h1ffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XConverter_4(
  input         io_in_clk,
  input         io_out_clk,
  input         io_rstn,
  input         io_in_valid,
  input  [31:0] io_in_bits_vaddr_high,
  input  [31:0] io_in_bits_vaddr_low,
  input  [31:0] io_in_bits_paddr_high,
  input  [31:0] io_in_bits_paddr_low,
  input         io_in_bits_is_base,
  output        io_out_valid,
  output [31:0] io_out_bits_vaddr_high,
  output [31:0] io_out_bits_vaddr_low,
  output [31:0] io_out_bits_paddr_high,
  output [31:0] io_out_bits_paddr_low,
  output        io_out_bits_is_base
);
  wire  fifo_io_m_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_s_clk; // @[XConverter.scala 97:34]
  wire  fifo_io_reset_n; // @[XConverter.scala 97:34]
  wire [135:0] fifo_io_in_data; // @[XConverter.scala 97:34]
  wire  fifo_io_in_valid; // @[XConverter.scala 97:34]
  wire [135:0] fifo_io_out_data; // @[XConverter.scala 97:34]
  wire  fifo_io_out_valid; // @[XConverter.scala 97:34]
  wire [128:0] _fifo_io_in_data_T = {io_in_bits_vaddr_high,io_in_bits_vaddr_low,io_in_bits_paddr_high,
    io_in_bits_paddr_low,io_in_bits_is_base}; // @[XConverter.scala 103:63]
  SV_STREAM_FIFO_4 fifo ( // @[XConverter.scala 97:34]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid)
  );
  assign io_out_valid = fifo_io_out_valid; // @[XConverter.scala 108:41]
  assign io_out_bits_vaddr_high = fifo_io_out_data[128:97]; // @[XConverter.scala 107:77]
  assign io_out_bits_vaddr_low = fifo_io_out_data[96:65]; // @[XConverter.scala 107:77]
  assign io_out_bits_paddr_high = fifo_io_out_data[64:33]; // @[XConverter.scala 107:77]
  assign io_out_bits_paddr_low = fifo_io_out_data[32:1]; // @[XConverter.scala 107:77]
  assign io_out_bits_is_base = fifo_io_out_data[0]; // @[XConverter.scala 107:77]
  assign fifo_io_m_clk = io_out_clk; // @[XConverter.scala 100:41]
  assign fifo_io_s_clk = io_in_clk; // @[XConverter.scala 99:41]
  assign fifo_io_reset_n = io_rstn; // @[XConverter.scala 101:41]
  assign fifo_io_in_data = {{7'd0}, _fifo_io_in_data_T}; // @[XConverter.scala 103:63]
  assign fifo_io_in_valid = io_in_valid; // @[XConverter.scala 104:41]
endmodule
module RegSlice(
  input         clock,
  input         reset,
  output        io_upStream_ready,
  input         io_upStream_valid,
  input  [31:0] io_upStream_bits_data,
  input         io_downStream_ready,
  output        io_downStream_valid,
  output [31:0] io_downStream_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  fwd_valid; // @[RegSlices.scala 112:34]
  reg [31:0] fwd_data_data; // @[RegSlices.scala 113:30]
  wire  fwd_ready_s = ~fwd_valid | io_downStream_ready; // @[RegSlices.scala 115:35]
  reg  bwd_ready; // @[RegSlices.scala 123:34]
  reg [31:0] bwd_data_data; // @[RegSlices.scala 124:30]
  wire  _fwd_valid_T = io_downStream_ready ? 1'h0 : fwd_valid; // @[RegSlices.scala 121:53]
  wire  bwd_valid_s = ~bwd_ready | io_upStream_valid; // @[RegSlices.scala 126:39]
  wire  _bwd_ready_T = io_upStream_valid ? 1'h0 : bwd_ready; // @[RegSlices.scala 132:53]
  assign io_upStream_ready = bwd_ready; // @[RegSlices.scala 107:31 RegSlices.scala 128:25]
  assign io_downStream_valid = fwd_valid; // @[RegSlices.scala 109:31 RegSlices.scala 116:21]
  assign io_downStream_bits_data = fwd_data_data; // @[RegSlices.scala 108:31 RegSlices.scala 117:25]
  always @(posedge clock) begin
    if (reset) begin // @[RegSlices.scala 112:34]
      fwd_valid <= 1'h0; // @[RegSlices.scala 112:34]
    end else begin
      fwd_valid <= bwd_valid_s | _fwd_valid_T; // @[RegSlices.scala 121:25]
    end
    if (fwd_ready_s) begin // @[RegSlices.scala 119:31]
      if (bwd_ready) begin // @[RegSlices.scala 127:31]
        fwd_data_data <= io_upStream_bits_data;
      end else begin
        fwd_data_data <= bwd_data_data;
      end
    end
    bwd_ready <= reset | (fwd_ready_s | _bwd_ready_T); // @[RegSlices.scala 123:34 RegSlices.scala 123:34 RegSlices.scala 132:25]
    if (bwd_ready) begin // @[RegSlices.scala 130:31]
      bwd_data_data <= io_upStream_bits_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fwd_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  fwd_data_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  bwd_ready = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  bwd_data_data = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PoorAXIL2Reg(
  input         clock,
  input         reset,
  output        io_axi_aw_ready,
  input         io_axi_aw_valid,
  input  [31:0] io_axi_aw_bits_addr,
  output        io_axi_ar_ready,
  input         io_axi_ar_valid,
  input  [31:0] io_axi_ar_bits_addr,
  output        io_axi_w_ready,
  input         io_axi_w_valid,
  input  [31:0] io_axi_w_bits_data,
  input         io_axi_r_ready,
  output        io_axi_r_valid,
  output [31:0] io_axi_r_bits_data,
  output [31:0] io_reg_control_8,
  output [31:0] io_reg_control_9,
  output [31:0] io_reg_control_10,
  output [31:0] io_reg_control_11,
  output [31:0] io_reg_control_12,
  output [31:0] io_reg_control_13,
  output [31:0] io_reg_control_20,
  output [31:0] io_reg_control_50,
  output [31:0] io_reg_control_51,
  output [31:0] io_reg_control_52,
  output [31:0] io_reg_control_53,
  output [31:0] io_reg_control_54,
  output [31:0] io_reg_control_55,
  output [31:0] io_reg_control_56,
  output [31:0] io_reg_control_57,
  output [31:0] io_reg_control_58,
  output [31:0] io_reg_control_59,
  output [31:0] io_reg_control_70,
  output [31:0] io_reg_control_71,
  output [31:0] io_reg_control_72,
  output [31:0] io_reg_control_73,
  output [31:0] io_reg_control_74,
  output [31:0] io_reg_control_75,
  output [31:0] io_reg_control_76,
  output [31:0] io_reg_control_77,
  output [31:0] io_reg_control_78,
  output [31:0] io_reg_control_79,
  output [31:0] io_reg_control_80,
  output [31:0] io_reg_control_91,
  output [31:0] io_reg_control_92,
  output [31:0] io_reg_control_93,
  output [31:0] io_reg_control_94,
  input  [31:0] io_reg_status_40,
  input  [31:0] io_reg_status_51,
  input  [31:0] io_reg_status_52,
  input  [31:0] io_reg_status_61,
  input  [31:0] io_reg_status_71,
  input  [31:0] io_reg_status_72,
  input  [31:0] io_reg_status_75,
  input  [31:0] io_reg_status_76,
  input  [31:0] io_reg_status_77,
  input  [31:0] io_reg_status_78,
  input  [31:0] io_reg_status_79,
  input  [31:0] io_reg_status_81
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
`endif // RANDOMIZE_REG_INIT
  wire  r_delay_clock; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_reset; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_io_upStream_ready; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_io_upStream_valid; // @[PoorAXIL2Reg.scala 38:33]
  wire [31:0] r_delay_io_upStream_bits_data; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_io_downStream_ready; // @[PoorAXIL2Reg.scala 38:33]
  wire  r_delay_io_downStream_valid; // @[PoorAXIL2Reg.scala 38:33]
  wire [31:0] r_delay_io_downStream_bits_data; // @[PoorAXIL2Reg.scala 38:33]
  reg [31:0] reg_control_8; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_9; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_10; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_11; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_12; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_13; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_20; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_50; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_51; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_52; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_53; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_54; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_55; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_56; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_57; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_58; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_59; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_70; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_71; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_72; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_73; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_74; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_75; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_76; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_77; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_78; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_79; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_80; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_91; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_92; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_93; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_control_94; // @[PoorAXIL2Reg.scala 17:30]
  reg [31:0] reg_status_40; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_51; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_52; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_61; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_71; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_72; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_75; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_76; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_77; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_78; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_79; // @[PoorAXIL2Reg.scala 19:29]
  reg [31:0] reg_status_81; // @[PoorAXIL2Reg.scala 19:29]
  reg  s_rd; // @[PoorAXIL2Reg.scala 30:27]
  reg  s_wr; // @[PoorAXIL2Reg.scala 31:27]
  reg [31:0] r_addr; // @[PoorAXIL2Reg.scala 41:25]
  reg [31:0] w_addr; // @[PoorAXIL2Reg.scala 42:25]
  wire  _io_axi_ar_ready_T = ~s_rd; // @[PoorAXIL2Reg.scala 44:74]
  wire [31:0] _GEN_40 = 9'h28 == r_addr[8:0] ? reg_status_40 : 32'h0; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_41 = 9'h29 == r_addr[8:0] ? 32'h0 : _GEN_40; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_42 = 9'h2a == r_addr[8:0] ? 32'h0 : _GEN_41; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_43 = 9'h2b == r_addr[8:0] ? 32'h0 : _GEN_42; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_44 = 9'h2c == r_addr[8:0] ? 32'h0 : _GEN_43; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_45 = 9'h2d == r_addr[8:0] ? 32'h0 : _GEN_44; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_46 = 9'h2e == r_addr[8:0] ? 32'h0 : _GEN_45; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_47 = 9'h2f == r_addr[8:0] ? 32'h0 : _GEN_46; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_48 = 9'h30 == r_addr[8:0] ? 32'h0 : _GEN_47; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_49 = 9'h31 == r_addr[8:0] ? 32'h0 : _GEN_48; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_50 = 9'h32 == r_addr[8:0] ? 32'h0 : _GEN_49; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_51 = 9'h33 == r_addr[8:0] ? reg_status_51 : _GEN_50; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_52 = 9'h34 == r_addr[8:0] ? reg_status_52 : _GEN_51; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_53 = 9'h35 == r_addr[8:0] ? 32'h0 : _GEN_52; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_54 = 9'h36 == r_addr[8:0] ? 32'h0 : _GEN_53; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_55 = 9'h37 == r_addr[8:0] ? 32'h0 : _GEN_54; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_56 = 9'h38 == r_addr[8:0] ? 32'h0 : _GEN_55; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_57 = 9'h39 == r_addr[8:0] ? 32'h0 : _GEN_56; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_58 = 9'h3a == r_addr[8:0] ? 32'h0 : _GEN_57; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_59 = 9'h3b == r_addr[8:0] ? 32'h0 : _GEN_58; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_60 = 9'h3c == r_addr[8:0] ? 32'h0 : _GEN_59; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_61 = 9'h3d == r_addr[8:0] ? reg_status_61 : _GEN_60; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_62 = 9'h3e == r_addr[8:0] ? 32'h0 : _GEN_61; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_63 = 9'h3f == r_addr[8:0] ? 32'h0 : _GEN_62; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_64 = 9'h40 == r_addr[8:0] ? 32'h0 : _GEN_63; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_65 = 9'h41 == r_addr[8:0] ? 32'h0 : _GEN_64; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_66 = 9'h42 == r_addr[8:0] ? 32'h0 : _GEN_65; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_67 = 9'h43 == r_addr[8:0] ? 32'h0 : _GEN_66; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_68 = 9'h44 == r_addr[8:0] ? 32'h0 : _GEN_67; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_69 = 9'h45 == r_addr[8:0] ? 32'h0 : _GEN_68; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_70 = 9'h46 == r_addr[8:0] ? 32'h0 : _GEN_69; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_71 = 9'h47 == r_addr[8:0] ? reg_status_71 : _GEN_70; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_72 = 9'h48 == r_addr[8:0] ? reg_status_72 : _GEN_71; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_73 = 9'h49 == r_addr[8:0] ? 32'h0 : _GEN_72; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_74 = 9'h4a == r_addr[8:0] ? 32'h0 : _GEN_73; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_75 = 9'h4b == r_addr[8:0] ? reg_status_75 : _GEN_74; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_76 = 9'h4c == r_addr[8:0] ? reg_status_76 : _GEN_75; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_77 = 9'h4d == r_addr[8:0] ? reg_status_77 : _GEN_76; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_78 = 9'h4e == r_addr[8:0] ? reg_status_78 : _GEN_77; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_79 = 9'h4f == r_addr[8:0] ? reg_status_79 : _GEN_78; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_80 = 9'h50 == r_addr[8:0] ? 32'h0 : _GEN_79; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_81 = 9'h51 == r_addr[8:0] ? reg_status_81 : _GEN_80; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_82 = 9'h52 == r_addr[8:0] ? 32'h0 : _GEN_81; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_83 = 9'h53 == r_addr[8:0] ? 32'h0 : _GEN_82; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_84 = 9'h54 == r_addr[8:0] ? 32'h0 : _GEN_83; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_85 = 9'h55 == r_addr[8:0] ? 32'h0 : _GEN_84; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_86 = 9'h56 == r_addr[8:0] ? 32'h0 : _GEN_85; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_87 = 9'h57 == r_addr[8:0] ? 32'h0 : _GEN_86; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_88 = 9'h58 == r_addr[8:0] ? 32'h0 : _GEN_87; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_89 = 9'h59 == r_addr[8:0] ? 32'h0 : _GEN_88; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_90 = 9'h5a == r_addr[8:0] ? 32'h0 : _GEN_89; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_91 = 9'h5b == r_addr[8:0] ? 32'h0 : _GEN_90; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_92 = 9'h5c == r_addr[8:0] ? 32'h0 : _GEN_91; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_93 = 9'h5d == r_addr[8:0] ? 32'h0 : _GEN_92; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_94 = 9'h5e == r_addr[8:0] ? 32'h0 : _GEN_93; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_95 = 9'h5f == r_addr[8:0] ? 32'h0 : _GEN_94; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_96 = 9'h60 == r_addr[8:0] ? 32'h0 : _GEN_95; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_97 = 9'h61 == r_addr[8:0] ? 32'h0 : _GEN_96; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_98 = 9'h62 == r_addr[8:0] ? 32'h0 : _GEN_97; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_99 = 9'h63 == r_addr[8:0] ? 32'h0 : _GEN_98; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_100 = 9'h64 == r_addr[8:0] ? 32'h0 : _GEN_99; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_101 = 9'h65 == r_addr[8:0] ? 32'h0 : _GEN_100; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_102 = 9'h66 == r_addr[8:0] ? 32'h0 : _GEN_101; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_103 = 9'h67 == r_addr[8:0] ? 32'h0 : _GEN_102; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_104 = 9'h68 == r_addr[8:0] ? 32'h0 : _GEN_103; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_105 = 9'h69 == r_addr[8:0] ? 32'h0 : _GEN_104; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_106 = 9'h6a == r_addr[8:0] ? 32'h0 : _GEN_105; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_107 = 9'h6b == r_addr[8:0] ? 32'h0 : _GEN_106; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_108 = 9'h6c == r_addr[8:0] ? 32'h0 : _GEN_107; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_109 = 9'h6d == r_addr[8:0] ? 32'h0 : _GEN_108; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_110 = 9'h6e == r_addr[8:0] ? 32'h0 : _GEN_109; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_111 = 9'h6f == r_addr[8:0] ? 32'h0 : _GEN_110; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_112 = 9'h70 == r_addr[8:0] ? 32'h0 : _GEN_111; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_113 = 9'h71 == r_addr[8:0] ? 32'h0 : _GEN_112; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_114 = 9'h72 == r_addr[8:0] ? 32'h0 : _GEN_113; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_115 = 9'h73 == r_addr[8:0] ? 32'h0 : _GEN_114; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_116 = 9'h74 == r_addr[8:0] ? 32'h0 : _GEN_115; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_117 = 9'h75 == r_addr[8:0] ? 32'h0 : _GEN_116; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_118 = 9'h76 == r_addr[8:0] ? 32'h0 : _GEN_117; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_119 = 9'h77 == r_addr[8:0] ? 32'h0 : _GEN_118; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_120 = 9'h78 == r_addr[8:0] ? 32'h0 : _GEN_119; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_121 = 9'h79 == r_addr[8:0] ? 32'h0 : _GEN_120; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_122 = 9'h7a == r_addr[8:0] ? 32'h0 : _GEN_121; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_123 = 9'h7b == r_addr[8:0] ? 32'h0 : _GEN_122; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_124 = 9'h7c == r_addr[8:0] ? 32'h0 : _GEN_123; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_125 = 9'h7d == r_addr[8:0] ? 32'h0 : _GEN_124; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_126 = 9'h7e == r_addr[8:0] ? 32'h0 : _GEN_125; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_127 = 9'h7f == r_addr[8:0] ? 32'h0 : _GEN_126; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_128 = 9'h80 == r_addr[8:0] ? 32'h0 : _GEN_127; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_129 = 9'h81 == r_addr[8:0] ? 32'h0 : _GEN_128; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_130 = 9'h82 == r_addr[8:0] ? 32'h0 : _GEN_129; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_131 = 9'h83 == r_addr[8:0] ? 32'h0 : _GEN_130; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_132 = 9'h84 == r_addr[8:0] ? 32'h0 : _GEN_131; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_133 = 9'h85 == r_addr[8:0] ? 32'h0 : _GEN_132; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_134 = 9'h86 == r_addr[8:0] ? 32'h0 : _GEN_133; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_135 = 9'h87 == r_addr[8:0] ? 32'h0 : _GEN_134; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_136 = 9'h88 == r_addr[8:0] ? 32'h0 : _GEN_135; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_137 = 9'h89 == r_addr[8:0] ? 32'h0 : _GEN_136; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_138 = 9'h8a == r_addr[8:0] ? 32'h0 : _GEN_137; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_139 = 9'h8b == r_addr[8:0] ? 32'h0 : _GEN_138; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_140 = 9'h8c == r_addr[8:0] ? 32'h0 : _GEN_139; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_141 = 9'h8d == r_addr[8:0] ? 32'h0 : _GEN_140; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_142 = 9'h8e == r_addr[8:0] ? 32'h0 : _GEN_141; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_143 = 9'h8f == r_addr[8:0] ? 32'h0 : _GEN_142; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_144 = 9'h90 == r_addr[8:0] ? 32'h0 : _GEN_143; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_145 = 9'h91 == r_addr[8:0] ? 32'h0 : _GEN_144; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_146 = 9'h92 == r_addr[8:0] ? 32'h0 : _GEN_145; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_147 = 9'h93 == r_addr[8:0] ? 32'h0 : _GEN_146; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_148 = 9'h94 == r_addr[8:0] ? 32'h0 : _GEN_147; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_149 = 9'h95 == r_addr[8:0] ? 32'h0 : _GEN_148; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_150 = 9'h96 == r_addr[8:0] ? 32'h0 : _GEN_149; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_151 = 9'h97 == r_addr[8:0] ? 32'h0 : _GEN_150; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_152 = 9'h98 == r_addr[8:0] ? 32'h0 : _GEN_151; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_153 = 9'h99 == r_addr[8:0] ? 32'h0 : _GEN_152; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_154 = 9'h9a == r_addr[8:0] ? 32'h0 : _GEN_153; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_155 = 9'h9b == r_addr[8:0] ? 32'h0 : _GEN_154; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_156 = 9'h9c == r_addr[8:0] ? 32'h0 : _GEN_155; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_157 = 9'h9d == r_addr[8:0] ? 32'h0 : _GEN_156; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_158 = 9'h9e == r_addr[8:0] ? 32'h0 : _GEN_157; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_159 = 9'h9f == r_addr[8:0] ? 32'h0 : _GEN_158; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_160 = 9'ha0 == r_addr[8:0] ? 32'h0 : _GEN_159; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_161 = 9'ha1 == r_addr[8:0] ? 32'h0 : _GEN_160; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_162 = 9'ha2 == r_addr[8:0] ? 32'h0 : _GEN_161; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_163 = 9'ha3 == r_addr[8:0] ? 32'h0 : _GEN_162; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_164 = 9'ha4 == r_addr[8:0] ? 32'h0 : _GEN_163; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_165 = 9'ha5 == r_addr[8:0] ? 32'h0 : _GEN_164; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_166 = 9'ha6 == r_addr[8:0] ? 32'h0 : _GEN_165; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_167 = 9'ha7 == r_addr[8:0] ? 32'h0 : _GEN_166; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_168 = 9'ha8 == r_addr[8:0] ? 32'h0 : _GEN_167; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_169 = 9'ha9 == r_addr[8:0] ? 32'h0 : _GEN_168; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_170 = 9'haa == r_addr[8:0] ? 32'h0 : _GEN_169; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_171 = 9'hab == r_addr[8:0] ? 32'h0 : _GEN_170; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_172 = 9'hac == r_addr[8:0] ? 32'h0 : _GEN_171; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_173 = 9'had == r_addr[8:0] ? 32'h0 : _GEN_172; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_174 = 9'hae == r_addr[8:0] ? 32'h0 : _GEN_173; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_175 = 9'haf == r_addr[8:0] ? 32'h0 : _GEN_174; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_176 = 9'hb0 == r_addr[8:0] ? 32'h0 : _GEN_175; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_177 = 9'hb1 == r_addr[8:0] ? 32'h0 : _GEN_176; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_178 = 9'hb2 == r_addr[8:0] ? 32'h0 : _GEN_177; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_179 = 9'hb3 == r_addr[8:0] ? 32'h0 : _GEN_178; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_180 = 9'hb4 == r_addr[8:0] ? 32'h0 : _GEN_179; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_181 = 9'hb5 == r_addr[8:0] ? 32'h0 : _GEN_180; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_182 = 9'hb6 == r_addr[8:0] ? 32'h0 : _GEN_181; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_183 = 9'hb7 == r_addr[8:0] ? 32'h0 : _GEN_182; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_184 = 9'hb8 == r_addr[8:0] ? 32'h0 : _GEN_183; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_185 = 9'hb9 == r_addr[8:0] ? 32'h0 : _GEN_184; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_186 = 9'hba == r_addr[8:0] ? 32'h0 : _GEN_185; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_187 = 9'hbb == r_addr[8:0] ? 32'h0 : _GEN_186; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_188 = 9'hbc == r_addr[8:0] ? 32'h0 : _GEN_187; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_189 = 9'hbd == r_addr[8:0] ? 32'h0 : _GEN_188; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_190 = 9'hbe == r_addr[8:0] ? 32'h0 : _GEN_189; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_191 = 9'hbf == r_addr[8:0] ? 32'h0 : _GEN_190; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_192 = 9'hc0 == r_addr[8:0] ? 32'h0 : _GEN_191; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_193 = 9'hc1 == r_addr[8:0] ? 32'h0 : _GEN_192; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_194 = 9'hc2 == r_addr[8:0] ? 32'h0 : _GEN_193; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_195 = 9'hc3 == r_addr[8:0] ? 32'h0 : _GEN_194; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_196 = 9'hc4 == r_addr[8:0] ? 32'h0 : _GEN_195; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_197 = 9'hc5 == r_addr[8:0] ? 32'h0 : _GEN_196; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_198 = 9'hc6 == r_addr[8:0] ? 32'h0 : _GEN_197; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_199 = 9'hc7 == r_addr[8:0] ? 32'h0 : _GEN_198; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_200 = 9'hc8 == r_addr[8:0] ? 32'h0 : _GEN_199; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_201 = 9'hc9 == r_addr[8:0] ? 32'h0 : _GEN_200; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_202 = 9'hca == r_addr[8:0] ? 32'h0 : _GEN_201; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_203 = 9'hcb == r_addr[8:0] ? 32'h0 : _GEN_202; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_204 = 9'hcc == r_addr[8:0] ? 32'h0 : _GEN_203; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_205 = 9'hcd == r_addr[8:0] ? 32'h0 : _GEN_204; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_206 = 9'hce == r_addr[8:0] ? 32'h0 : _GEN_205; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_207 = 9'hcf == r_addr[8:0] ? 32'h0 : _GEN_206; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_208 = 9'hd0 == r_addr[8:0] ? 32'h0 : _GEN_207; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_209 = 9'hd1 == r_addr[8:0] ? 32'h0 : _GEN_208; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_210 = 9'hd2 == r_addr[8:0] ? 32'h0 : _GEN_209; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_211 = 9'hd3 == r_addr[8:0] ? 32'h0 : _GEN_210; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_212 = 9'hd4 == r_addr[8:0] ? 32'h0 : _GEN_211; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_213 = 9'hd5 == r_addr[8:0] ? 32'h0 : _GEN_212; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_214 = 9'hd6 == r_addr[8:0] ? 32'h0 : _GEN_213; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_215 = 9'hd7 == r_addr[8:0] ? 32'h0 : _GEN_214; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_216 = 9'hd8 == r_addr[8:0] ? 32'h0 : _GEN_215; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_217 = 9'hd9 == r_addr[8:0] ? 32'h0 : _GEN_216; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_218 = 9'hda == r_addr[8:0] ? 32'h0 : _GEN_217; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_219 = 9'hdb == r_addr[8:0] ? 32'h0 : _GEN_218; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_220 = 9'hdc == r_addr[8:0] ? 32'h0 : _GEN_219; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_221 = 9'hdd == r_addr[8:0] ? 32'h0 : _GEN_220; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_222 = 9'hde == r_addr[8:0] ? 32'h0 : _GEN_221; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_223 = 9'hdf == r_addr[8:0] ? 32'h0 : _GEN_222; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_224 = 9'he0 == r_addr[8:0] ? 32'h0 : _GEN_223; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_225 = 9'he1 == r_addr[8:0] ? 32'h0 : _GEN_224; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_226 = 9'he2 == r_addr[8:0] ? 32'h0 : _GEN_225; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_227 = 9'he3 == r_addr[8:0] ? 32'h0 : _GEN_226; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_228 = 9'he4 == r_addr[8:0] ? 32'h0 : _GEN_227; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_229 = 9'he5 == r_addr[8:0] ? 32'h0 : _GEN_228; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_230 = 9'he6 == r_addr[8:0] ? 32'h0 : _GEN_229; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_231 = 9'he7 == r_addr[8:0] ? 32'h0 : _GEN_230; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_232 = 9'he8 == r_addr[8:0] ? 32'h0 : _GEN_231; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_233 = 9'he9 == r_addr[8:0] ? 32'h0 : _GEN_232; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_234 = 9'hea == r_addr[8:0] ? 32'h0 : _GEN_233; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_235 = 9'heb == r_addr[8:0] ? 32'h0 : _GEN_234; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_236 = 9'hec == r_addr[8:0] ? 32'h0 : _GEN_235; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_237 = 9'hed == r_addr[8:0] ? 32'h0 : _GEN_236; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_238 = 9'hee == r_addr[8:0] ? 32'h0 : _GEN_237; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_239 = 9'hef == r_addr[8:0] ? 32'h0 : _GEN_238; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_240 = 9'hf0 == r_addr[8:0] ? 32'h0 : _GEN_239; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_241 = 9'hf1 == r_addr[8:0] ? 32'h0 : _GEN_240; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_242 = 9'hf2 == r_addr[8:0] ? 32'h0 : _GEN_241; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_243 = 9'hf3 == r_addr[8:0] ? 32'h0 : _GEN_242; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_244 = 9'hf4 == r_addr[8:0] ? 32'h0 : _GEN_243; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_245 = 9'hf5 == r_addr[8:0] ? 32'h0 : _GEN_244; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_246 = 9'hf6 == r_addr[8:0] ? 32'h0 : _GEN_245; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_247 = 9'hf7 == r_addr[8:0] ? 32'h0 : _GEN_246; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_248 = 9'hf8 == r_addr[8:0] ? 32'h0 : _GEN_247; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_249 = 9'hf9 == r_addr[8:0] ? 32'h0 : _GEN_248; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_250 = 9'hfa == r_addr[8:0] ? 32'h0 : _GEN_249; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_251 = 9'hfb == r_addr[8:0] ? 32'h0 : _GEN_250; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_252 = 9'hfc == r_addr[8:0] ? 32'h0 : _GEN_251; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_253 = 9'hfd == r_addr[8:0] ? 32'h0 : _GEN_252; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_254 = 9'hfe == r_addr[8:0] ? 32'h0 : _GEN_253; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_255 = 9'hff == r_addr[8:0] ? 32'h0 : _GEN_254; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_256 = 9'h100 == r_addr[8:0] ? 32'h0 : _GEN_255; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_257 = 9'h101 == r_addr[8:0] ? 32'h0 : _GEN_256; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_258 = 9'h102 == r_addr[8:0] ? 32'h0 : _GEN_257; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_259 = 9'h103 == r_addr[8:0] ? 32'h0 : _GEN_258; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_260 = 9'h104 == r_addr[8:0] ? 32'h0 : _GEN_259; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_261 = 9'h105 == r_addr[8:0] ? 32'h0 : _GEN_260; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_262 = 9'h106 == r_addr[8:0] ? 32'h0 : _GEN_261; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_263 = 9'h107 == r_addr[8:0] ? 32'h0 : _GEN_262; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_264 = 9'h108 == r_addr[8:0] ? 32'h0 : _GEN_263; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_265 = 9'h109 == r_addr[8:0] ? 32'h0 : _GEN_264; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_266 = 9'h10a == r_addr[8:0] ? 32'h0 : _GEN_265; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_267 = 9'h10b == r_addr[8:0] ? 32'h0 : _GEN_266; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_268 = 9'h10c == r_addr[8:0] ? 32'h0 : _GEN_267; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_269 = 9'h10d == r_addr[8:0] ? 32'h0 : _GEN_268; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_270 = 9'h10e == r_addr[8:0] ? 32'h0 : _GEN_269; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_271 = 9'h10f == r_addr[8:0] ? 32'h0 : _GEN_270; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_272 = 9'h110 == r_addr[8:0] ? 32'h0 : _GEN_271; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_273 = 9'h111 == r_addr[8:0] ? 32'h0 : _GEN_272; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_274 = 9'h112 == r_addr[8:0] ? 32'h0 : _GEN_273; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_275 = 9'h113 == r_addr[8:0] ? 32'h0 : _GEN_274; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_276 = 9'h114 == r_addr[8:0] ? 32'h0 : _GEN_275; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_277 = 9'h115 == r_addr[8:0] ? 32'h0 : _GEN_276; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_278 = 9'h116 == r_addr[8:0] ? 32'h0 : _GEN_277; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_279 = 9'h117 == r_addr[8:0] ? 32'h0 : _GEN_278; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_280 = 9'h118 == r_addr[8:0] ? 32'h0 : _GEN_279; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_281 = 9'h119 == r_addr[8:0] ? 32'h0 : _GEN_280; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_282 = 9'h11a == r_addr[8:0] ? 32'h0 : _GEN_281; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_283 = 9'h11b == r_addr[8:0] ? 32'h0 : _GEN_282; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_284 = 9'h11c == r_addr[8:0] ? 32'h0 : _GEN_283; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_285 = 9'h11d == r_addr[8:0] ? 32'h0 : _GEN_284; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_286 = 9'h11e == r_addr[8:0] ? 32'h0 : _GEN_285; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_287 = 9'h11f == r_addr[8:0] ? 32'h0 : _GEN_286; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_288 = 9'h120 == r_addr[8:0] ? 32'h0 : _GEN_287; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_289 = 9'h121 == r_addr[8:0] ? 32'h0 : _GEN_288; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_290 = 9'h122 == r_addr[8:0] ? 32'h0 : _GEN_289; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_291 = 9'h123 == r_addr[8:0] ? 32'h0 : _GEN_290; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_292 = 9'h124 == r_addr[8:0] ? 32'h0 : _GEN_291; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_293 = 9'h125 == r_addr[8:0] ? 32'h0 : _GEN_292; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_294 = 9'h126 == r_addr[8:0] ? 32'h0 : _GEN_293; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_295 = 9'h127 == r_addr[8:0] ? 32'h0 : _GEN_294; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_296 = 9'h128 == r_addr[8:0] ? 32'h0 : _GEN_295; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_297 = 9'h129 == r_addr[8:0] ? 32'h0 : _GEN_296; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_298 = 9'h12a == r_addr[8:0] ? 32'h0 : _GEN_297; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_299 = 9'h12b == r_addr[8:0] ? 32'h0 : _GEN_298; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_300 = 9'h12c == r_addr[8:0] ? 32'h0 : _GEN_299; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_301 = 9'h12d == r_addr[8:0] ? 32'h0 : _GEN_300; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_302 = 9'h12e == r_addr[8:0] ? 32'h0 : _GEN_301; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_303 = 9'h12f == r_addr[8:0] ? 32'h0 : _GEN_302; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_304 = 9'h130 == r_addr[8:0] ? 32'h0 : _GEN_303; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_305 = 9'h131 == r_addr[8:0] ? 32'h0 : _GEN_304; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_306 = 9'h132 == r_addr[8:0] ? 32'h0 : _GEN_305; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_307 = 9'h133 == r_addr[8:0] ? 32'h0 : _GEN_306; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_308 = 9'h134 == r_addr[8:0] ? 32'h0 : _GEN_307; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_309 = 9'h135 == r_addr[8:0] ? 32'h0 : _GEN_308; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_310 = 9'h136 == r_addr[8:0] ? 32'h0 : _GEN_309; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_311 = 9'h137 == r_addr[8:0] ? 32'h0 : _GEN_310; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_312 = 9'h138 == r_addr[8:0] ? 32'h0 : _GEN_311; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_313 = 9'h139 == r_addr[8:0] ? 32'h0 : _GEN_312; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_314 = 9'h13a == r_addr[8:0] ? 32'h0 : _GEN_313; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_315 = 9'h13b == r_addr[8:0] ? 32'h0 : _GEN_314; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_316 = 9'h13c == r_addr[8:0] ? 32'h0 : _GEN_315; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_317 = 9'h13d == r_addr[8:0] ? 32'h0 : _GEN_316; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_318 = 9'h13e == r_addr[8:0] ? 32'h0 : _GEN_317; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_319 = 9'h13f == r_addr[8:0] ? 32'h0 : _GEN_318; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_320 = 9'h140 == r_addr[8:0] ? 32'h0 : _GEN_319; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_321 = 9'h141 == r_addr[8:0] ? 32'h0 : _GEN_320; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_322 = 9'h142 == r_addr[8:0] ? 32'h0 : _GEN_321; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_323 = 9'h143 == r_addr[8:0] ? 32'h0 : _GEN_322; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_324 = 9'h144 == r_addr[8:0] ? 32'h0 : _GEN_323; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_325 = 9'h145 == r_addr[8:0] ? 32'h0 : _GEN_324; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_326 = 9'h146 == r_addr[8:0] ? 32'h0 : _GEN_325; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_327 = 9'h147 == r_addr[8:0] ? 32'h0 : _GEN_326; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_328 = 9'h148 == r_addr[8:0] ? 32'h0 : _GEN_327; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_329 = 9'h149 == r_addr[8:0] ? 32'h0 : _GEN_328; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_330 = 9'h14a == r_addr[8:0] ? 32'h0 : _GEN_329; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_331 = 9'h14b == r_addr[8:0] ? 32'h0 : _GEN_330; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_332 = 9'h14c == r_addr[8:0] ? 32'h0 : _GEN_331; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_333 = 9'h14d == r_addr[8:0] ? 32'h0 : _GEN_332; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_334 = 9'h14e == r_addr[8:0] ? 32'h0 : _GEN_333; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_335 = 9'h14f == r_addr[8:0] ? 32'h0 : _GEN_334; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_336 = 9'h150 == r_addr[8:0] ? 32'h0 : _GEN_335; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_337 = 9'h151 == r_addr[8:0] ? 32'h0 : _GEN_336; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_338 = 9'h152 == r_addr[8:0] ? 32'h0 : _GEN_337; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_339 = 9'h153 == r_addr[8:0] ? 32'h0 : _GEN_338; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_340 = 9'h154 == r_addr[8:0] ? 32'h0 : _GEN_339; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_341 = 9'h155 == r_addr[8:0] ? 32'h0 : _GEN_340; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_342 = 9'h156 == r_addr[8:0] ? 32'h0 : _GEN_341; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_343 = 9'h157 == r_addr[8:0] ? 32'h0 : _GEN_342; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_344 = 9'h158 == r_addr[8:0] ? 32'h0 : _GEN_343; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_345 = 9'h159 == r_addr[8:0] ? 32'h0 : _GEN_344; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_346 = 9'h15a == r_addr[8:0] ? 32'h0 : _GEN_345; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_347 = 9'h15b == r_addr[8:0] ? 32'h0 : _GEN_346; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_348 = 9'h15c == r_addr[8:0] ? 32'h0 : _GEN_347; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_349 = 9'h15d == r_addr[8:0] ? 32'h0 : _GEN_348; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_350 = 9'h15e == r_addr[8:0] ? 32'h0 : _GEN_349; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_351 = 9'h15f == r_addr[8:0] ? 32'h0 : _GEN_350; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_352 = 9'h160 == r_addr[8:0] ? 32'h0 : _GEN_351; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_353 = 9'h161 == r_addr[8:0] ? 32'h0 : _GEN_352; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_354 = 9'h162 == r_addr[8:0] ? 32'h0 : _GEN_353; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_355 = 9'h163 == r_addr[8:0] ? 32'h0 : _GEN_354; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_356 = 9'h164 == r_addr[8:0] ? 32'h0 : _GEN_355; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_357 = 9'h165 == r_addr[8:0] ? 32'h0 : _GEN_356; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_358 = 9'h166 == r_addr[8:0] ? 32'h0 : _GEN_357; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_359 = 9'h167 == r_addr[8:0] ? 32'h0 : _GEN_358; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_360 = 9'h168 == r_addr[8:0] ? 32'h0 : _GEN_359; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_361 = 9'h169 == r_addr[8:0] ? 32'h0 : _GEN_360; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_362 = 9'h16a == r_addr[8:0] ? 32'h0 : _GEN_361; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_363 = 9'h16b == r_addr[8:0] ? 32'h0 : _GEN_362; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_364 = 9'h16c == r_addr[8:0] ? 32'h0 : _GEN_363; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_365 = 9'h16d == r_addr[8:0] ? 32'h0 : _GEN_364; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_366 = 9'h16e == r_addr[8:0] ? 32'h0 : _GEN_365; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_367 = 9'h16f == r_addr[8:0] ? 32'h0 : _GEN_366; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_368 = 9'h170 == r_addr[8:0] ? 32'h0 : _GEN_367; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_369 = 9'h171 == r_addr[8:0] ? 32'h0 : _GEN_368; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_370 = 9'h172 == r_addr[8:0] ? 32'h0 : _GEN_369; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_371 = 9'h173 == r_addr[8:0] ? 32'h0 : _GEN_370; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_372 = 9'h174 == r_addr[8:0] ? 32'h0 : _GEN_371; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_373 = 9'h175 == r_addr[8:0] ? 32'h0 : _GEN_372; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_374 = 9'h176 == r_addr[8:0] ? 32'h0 : _GEN_373; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_375 = 9'h177 == r_addr[8:0] ? 32'h0 : _GEN_374; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_376 = 9'h178 == r_addr[8:0] ? 32'h0 : _GEN_375; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_377 = 9'h179 == r_addr[8:0] ? 32'h0 : _GEN_376; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_378 = 9'h17a == r_addr[8:0] ? 32'h0 : _GEN_377; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_379 = 9'h17b == r_addr[8:0] ? 32'h0 : _GEN_378; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_380 = 9'h17c == r_addr[8:0] ? 32'h0 : _GEN_379; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_381 = 9'h17d == r_addr[8:0] ? 32'h0 : _GEN_380; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_382 = 9'h17e == r_addr[8:0] ? 32'h0 : _GEN_381; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_383 = 9'h17f == r_addr[8:0] ? 32'h0 : _GEN_382; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_384 = 9'h180 == r_addr[8:0] ? 32'h0 : _GEN_383; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_385 = 9'h181 == r_addr[8:0] ? 32'h0 : _GEN_384; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_386 = 9'h182 == r_addr[8:0] ? 32'h0 : _GEN_385; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_387 = 9'h183 == r_addr[8:0] ? 32'h0 : _GEN_386; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_388 = 9'h184 == r_addr[8:0] ? 32'h0 : _GEN_387; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_389 = 9'h185 == r_addr[8:0] ? 32'h0 : _GEN_388; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_390 = 9'h186 == r_addr[8:0] ? 32'h0 : _GEN_389; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_391 = 9'h187 == r_addr[8:0] ? 32'h0 : _GEN_390; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_392 = 9'h188 == r_addr[8:0] ? 32'h0 : _GEN_391; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_393 = 9'h189 == r_addr[8:0] ? 32'h0 : _GEN_392; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_394 = 9'h18a == r_addr[8:0] ? 32'h0 : _GEN_393; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_395 = 9'h18b == r_addr[8:0] ? 32'h0 : _GEN_394; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_396 = 9'h18c == r_addr[8:0] ? 32'h0 : _GEN_395; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_397 = 9'h18d == r_addr[8:0] ? 32'h0 : _GEN_396; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_398 = 9'h18e == r_addr[8:0] ? 32'h0 : _GEN_397; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_399 = 9'h18f == r_addr[8:0] ? 32'h0 : _GEN_398; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_400 = 9'h190 == r_addr[8:0] ? 32'h0 : _GEN_399; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_401 = 9'h191 == r_addr[8:0] ? 32'h0 : _GEN_400; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_402 = 9'h192 == r_addr[8:0] ? 32'h0 : _GEN_401; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_403 = 9'h193 == r_addr[8:0] ? 32'h0 : _GEN_402; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_404 = 9'h194 == r_addr[8:0] ? 32'h0 : _GEN_403; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_405 = 9'h195 == r_addr[8:0] ? 32'h0 : _GEN_404; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_406 = 9'h196 == r_addr[8:0] ? 32'h0 : _GEN_405; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_407 = 9'h197 == r_addr[8:0] ? 32'h0 : _GEN_406; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_408 = 9'h198 == r_addr[8:0] ? 32'h0 : _GEN_407; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_409 = 9'h199 == r_addr[8:0] ? 32'h0 : _GEN_408; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_410 = 9'h19a == r_addr[8:0] ? 32'h0 : _GEN_409; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_411 = 9'h19b == r_addr[8:0] ? 32'h0 : _GEN_410; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_412 = 9'h19c == r_addr[8:0] ? 32'h0 : _GEN_411; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_413 = 9'h19d == r_addr[8:0] ? 32'h0 : _GEN_412; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_414 = 9'h19e == r_addr[8:0] ? 32'h0 : _GEN_413; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_415 = 9'h19f == r_addr[8:0] ? 32'h0 : _GEN_414; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_416 = 9'h1a0 == r_addr[8:0] ? 32'h0 : _GEN_415; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_417 = 9'h1a1 == r_addr[8:0] ? 32'h0 : _GEN_416; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_418 = 9'h1a2 == r_addr[8:0] ? 32'h0 : _GEN_417; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_419 = 9'h1a3 == r_addr[8:0] ? 32'h0 : _GEN_418; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_420 = 9'h1a4 == r_addr[8:0] ? 32'h0 : _GEN_419; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_421 = 9'h1a5 == r_addr[8:0] ? 32'h0 : _GEN_420; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_422 = 9'h1a6 == r_addr[8:0] ? 32'h0 : _GEN_421; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_423 = 9'h1a7 == r_addr[8:0] ? 32'h0 : _GEN_422; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_424 = 9'h1a8 == r_addr[8:0] ? 32'h0 : _GEN_423; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_425 = 9'h1a9 == r_addr[8:0] ? 32'h0 : _GEN_424; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_426 = 9'h1aa == r_addr[8:0] ? 32'h0 : _GEN_425; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_427 = 9'h1ab == r_addr[8:0] ? 32'h0 : _GEN_426; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_428 = 9'h1ac == r_addr[8:0] ? 32'h0 : _GEN_427; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_429 = 9'h1ad == r_addr[8:0] ? 32'h0 : _GEN_428; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_430 = 9'h1ae == r_addr[8:0] ? 32'h0 : _GEN_429; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_431 = 9'h1af == r_addr[8:0] ? 32'h0 : _GEN_430; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_432 = 9'h1b0 == r_addr[8:0] ? 32'h0 : _GEN_431; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_433 = 9'h1b1 == r_addr[8:0] ? 32'h0 : _GEN_432; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_434 = 9'h1b2 == r_addr[8:0] ? 32'h0 : _GEN_433; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_435 = 9'h1b3 == r_addr[8:0] ? 32'h0 : _GEN_434; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_436 = 9'h1b4 == r_addr[8:0] ? 32'h0 : _GEN_435; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_437 = 9'h1b5 == r_addr[8:0] ? 32'h0 : _GEN_436; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_438 = 9'h1b6 == r_addr[8:0] ? 32'h0 : _GEN_437; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_439 = 9'h1b7 == r_addr[8:0] ? 32'h0 : _GEN_438; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_440 = 9'h1b8 == r_addr[8:0] ? 32'h0 : _GEN_439; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_441 = 9'h1b9 == r_addr[8:0] ? 32'h0 : _GEN_440; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_442 = 9'h1ba == r_addr[8:0] ? 32'h0 : _GEN_441; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_443 = 9'h1bb == r_addr[8:0] ? 32'h0 : _GEN_442; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_444 = 9'h1bc == r_addr[8:0] ? 32'h0 : _GEN_443; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_445 = 9'h1bd == r_addr[8:0] ? 32'h0 : _GEN_444; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_446 = 9'h1be == r_addr[8:0] ? 32'h0 : _GEN_445; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_447 = 9'h1bf == r_addr[8:0] ? 32'h0 : _GEN_446; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_448 = 9'h1c0 == r_addr[8:0] ? 32'h0 : _GEN_447; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_449 = 9'h1c1 == r_addr[8:0] ? 32'h0 : _GEN_448; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_450 = 9'h1c2 == r_addr[8:0] ? 32'h0 : _GEN_449; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_451 = 9'h1c3 == r_addr[8:0] ? 32'h0 : _GEN_450; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_452 = 9'h1c4 == r_addr[8:0] ? 32'h0 : _GEN_451; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_453 = 9'h1c5 == r_addr[8:0] ? 32'h0 : _GEN_452; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_454 = 9'h1c6 == r_addr[8:0] ? 32'h0 : _GEN_453; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_455 = 9'h1c7 == r_addr[8:0] ? 32'h0 : _GEN_454; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_456 = 9'h1c8 == r_addr[8:0] ? 32'h0 : _GEN_455; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_457 = 9'h1c9 == r_addr[8:0] ? 32'h0 : _GEN_456; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_458 = 9'h1ca == r_addr[8:0] ? 32'h0 : _GEN_457; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_459 = 9'h1cb == r_addr[8:0] ? 32'h0 : _GEN_458; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_460 = 9'h1cc == r_addr[8:0] ? 32'h0 : _GEN_459; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_461 = 9'h1cd == r_addr[8:0] ? 32'h0 : _GEN_460; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_462 = 9'h1ce == r_addr[8:0] ? 32'h0 : _GEN_461; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_463 = 9'h1cf == r_addr[8:0] ? 32'h0 : _GEN_462; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_464 = 9'h1d0 == r_addr[8:0] ? 32'h0 : _GEN_463; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_465 = 9'h1d1 == r_addr[8:0] ? 32'h0 : _GEN_464; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_466 = 9'h1d2 == r_addr[8:0] ? 32'h0 : _GEN_465; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_467 = 9'h1d3 == r_addr[8:0] ? 32'h0 : _GEN_466; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_468 = 9'h1d4 == r_addr[8:0] ? 32'h0 : _GEN_467; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_469 = 9'h1d5 == r_addr[8:0] ? 32'h0 : _GEN_468; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_470 = 9'h1d6 == r_addr[8:0] ? 32'h0 : _GEN_469; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_471 = 9'h1d7 == r_addr[8:0] ? 32'h0 : _GEN_470; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_472 = 9'h1d8 == r_addr[8:0] ? 32'h0 : _GEN_471; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_473 = 9'h1d9 == r_addr[8:0] ? 32'h0 : _GEN_472; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_474 = 9'h1da == r_addr[8:0] ? 32'h0 : _GEN_473; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_475 = 9'h1db == r_addr[8:0] ? 32'h0 : _GEN_474; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_476 = 9'h1dc == r_addr[8:0] ? 32'h0 : _GEN_475; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_477 = 9'h1dd == r_addr[8:0] ? 32'h0 : _GEN_476; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_478 = 9'h1de == r_addr[8:0] ? 32'h0 : _GEN_477; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_479 = 9'h1df == r_addr[8:0] ? 32'h0 : _GEN_478; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_480 = 9'h1e0 == r_addr[8:0] ? 32'h0 : _GEN_479; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_481 = 9'h1e1 == r_addr[8:0] ? 32'h0 : _GEN_480; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_482 = 9'h1e2 == r_addr[8:0] ? 32'h0 : _GEN_481; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_483 = 9'h1e3 == r_addr[8:0] ? 32'h0 : _GEN_482; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_484 = 9'h1e4 == r_addr[8:0] ? 32'h0 : _GEN_483; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_485 = 9'h1e5 == r_addr[8:0] ? 32'h0 : _GEN_484; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_486 = 9'h1e6 == r_addr[8:0] ? 32'h0 : _GEN_485; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_487 = 9'h1e7 == r_addr[8:0] ? 32'h0 : _GEN_486; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_488 = 9'h1e8 == r_addr[8:0] ? 32'h0 : _GEN_487; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_489 = 9'h1e9 == r_addr[8:0] ? 32'h0 : _GEN_488; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_490 = 9'h1ea == r_addr[8:0] ? 32'h0 : _GEN_489; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_491 = 9'h1eb == r_addr[8:0] ? 32'h0 : _GEN_490; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_492 = 9'h1ec == r_addr[8:0] ? 32'h0 : _GEN_491; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_493 = 9'h1ed == r_addr[8:0] ? 32'h0 : _GEN_492; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_494 = 9'h1ee == r_addr[8:0] ? 32'h0 : _GEN_493; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_495 = 9'h1ef == r_addr[8:0] ? 32'h0 : _GEN_494; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_496 = 9'h1f0 == r_addr[8:0] ? 32'h0 : _GEN_495; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_497 = 9'h1f1 == r_addr[8:0] ? 32'h0 : _GEN_496; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_498 = 9'h1f2 == r_addr[8:0] ? 32'h0 : _GEN_497; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_499 = 9'h1f3 == r_addr[8:0] ? 32'h0 : _GEN_498; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_500 = 9'h1f4 == r_addr[8:0] ? 32'h0 : _GEN_499; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_501 = 9'h1f5 == r_addr[8:0] ? 32'h0 : _GEN_500; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_502 = 9'h1f6 == r_addr[8:0] ? 32'h0 : _GEN_501; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_503 = 9'h1f7 == r_addr[8:0] ? 32'h0 : _GEN_502; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_504 = 9'h1f8 == r_addr[8:0] ? 32'h0 : _GEN_503; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_505 = 9'h1f9 == r_addr[8:0] ? 32'h0 : _GEN_504; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_506 = 9'h1fa == r_addr[8:0] ? 32'h0 : _GEN_505; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_507 = 9'h1fb == r_addr[8:0] ? 32'h0 : _GEN_506; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_508 = 9'h1fc == r_addr[8:0] ? 32'h0 : _GEN_507; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_509 = 9'h1fd == r_addr[8:0] ? 32'h0 : _GEN_508; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire [31:0] _GEN_510 = 9'h1fe == r_addr[8:0] ? 32'h0 : _GEN_509; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  wire  _T_1 = io_axi_ar_ready & io_axi_ar_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _r_addr_T = {{2'd0}, io_axi_ar_bits_addr[31:2]}; // @[PoorAXIL2Reg.scala 51:73]
  wire  _GEN_513 = _T_1 | s_rd; // @[PoorAXIL2Reg.scala 50:40 PoorAXIL2Reg.scala 52:57 PoorAXIL2Reg.scala 30:27]
  wire  _T_3 = r_delay_io_upStream_ready & r_delay_io_upStream_valid; // @[Decoupled.scala 40:37]
  wire  _io_axi_aw_ready_T = ~s_wr; // @[PoorAXIL2Reg.scala 62:34]
  wire  _T_4 = io_axi_w_ready & io_axi_w_valid; // @[Decoupled.scala 40:37]
  wire  _T_7 = io_axi_aw_ready & io_axi_aw_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _w_addr_T = {{2'd0}, io_axi_aw_bits_addr[31:2]}; // @[PoorAXIL2Reg.scala 70:73]
  wire  _GEN_1543 = _T_7 | s_wr; // @[PoorAXIL2Reg.scala 69:40 PoorAXIL2Reg.scala 71:57 PoorAXIL2Reg.scala 31:27]
  RegSlice r_delay ( // @[PoorAXIL2Reg.scala 38:33]
    .clock(r_delay_clock),
    .reset(r_delay_reset),
    .io_upStream_ready(r_delay_io_upStream_ready),
    .io_upStream_valid(r_delay_io_upStream_valid),
    .io_upStream_bits_data(r_delay_io_upStream_bits_data),
    .io_downStream_ready(r_delay_io_downStream_ready),
    .io_downStream_valid(r_delay_io_downStream_valid),
    .io_downStream_bits_data(r_delay_io_downStream_bits_data)
  );
  assign io_axi_aw_ready = ~s_wr; // @[PoorAXIL2Reg.scala 62:34]
  assign io_axi_ar_ready = ~s_rd; // @[PoorAXIL2Reg.scala 44:74]
  assign io_axi_w_ready = s_wr; // @[PoorAXIL2Reg.scala 63:34]
  assign io_axi_r_valid = r_delay_io_downStream_valid; // @[PoorAXIL2Reg.scala 47:73]
  assign io_axi_r_bits_data = r_delay_io_downStream_bits_data; // @[PoorAXIL2Reg.scala 47:73]
  assign io_reg_control_8 = reg_control_8; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_9 = reg_control_9; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_10 = reg_control_10; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_11 = reg_control_11; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_12 = reg_control_12; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_13 = reg_control_13; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_20 = reg_control_20; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_50 = reg_control_50; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_51 = reg_control_51; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_52 = reg_control_52; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_53 = reg_control_53; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_54 = reg_control_54; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_55 = reg_control_55; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_56 = reg_control_56; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_57 = reg_control_57; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_58 = reg_control_58; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_59 = reg_control_59; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_70 = reg_control_70; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_71 = reg_control_71; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_72 = reg_control_72; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_73 = reg_control_73; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_74 = reg_control_74; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_75 = reg_control_75; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_76 = reg_control_76; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_77 = reg_control_77; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_78 = reg_control_78; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_79 = reg_control_79; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_80 = reg_control_80; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_91 = reg_control_91; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_92 = reg_control_92; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_93 = reg_control_93; // @[PoorAXIL2Reg.scala 23:57]
  assign io_reg_control_94 = reg_control_94; // @[PoorAXIL2Reg.scala 23:57]
  assign r_delay_clock = clock;
  assign r_delay_reset = reset;
  assign r_delay_io_upStream_valid = s_rd; // @[PoorAXIL2Reg.scala 45:58]
  assign r_delay_io_upStream_bits_data = 9'h1ff == r_addr[8:0] ? 32'h0 : _GEN_510; // @[PoorAXIL2Reg.scala 46:41 PoorAXIL2Reg.scala 46:41]
  assign r_delay_io_downStream_ready = io_axi_r_ready; // @[PoorAXIL2Reg.scala 47:73]
  always @(posedge clock) begin
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h8 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_8 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h9 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_9 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'ha == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_10 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'hb == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_11 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'hc == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_12 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'hd == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_13 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h14 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_20 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h32 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_50 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h33 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_51 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h34 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_52 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h35 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_53 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h36 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_54 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h37 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_55 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h38 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_56 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h39 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_57 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h3a == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_58 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h3b == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_59 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h46 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_70 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h47 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_71 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h48 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_72 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h49 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_73 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h4a == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_74 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h4b == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_75 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h4c == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_76 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h4d == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_77 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h4e == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_78 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h4f == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_79 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h50 == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_80 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h5b == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_91 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h5c == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_92 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h5d == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_93 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    if (_T_4) begin // @[PoorAXIL2Reg.scala 64:23]
      if (9'h5e == w_addr[8:0]) begin // @[PoorAXIL2Reg.scala 65:41]
        reg_control_94 <= io_axi_w_bits_data; // @[PoorAXIL2Reg.scala 65:41]
      end
    end
    reg_status_40 <= io_reg_status_40; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_51 <= io_reg_status_51; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_52 <= io_reg_status_52; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_61 <= io_reg_status_61; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_71 <= io_reg_status_71; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_72 <= io_reg_status_72; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_75 <= io_reg_status_75; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_76 <= io_reg_status_76; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_77 <= io_reg_status_77; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_78 <= io_reg_status_78; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_79 <= io_reg_status_79; // @[PoorAXIL2Reg.scala 22:57]
    reg_status_81 <= io_reg_status_81; // @[PoorAXIL2Reg.scala 22:57]
    if (reset) begin // @[PoorAXIL2Reg.scala 30:27]
      s_rd <= 1'h0; // @[PoorAXIL2Reg.scala 30:27]
    end else if (_io_axi_ar_ready_T) begin // @[Conditional.scala 40:58]
      s_rd <= _GEN_513;
    end else if (s_rd) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[PoorAXIL2Reg.scala 56:57]
        s_rd <= 1'h0; // @[PoorAXIL2Reg.scala 57:57]
      end
    end
    if (reset) begin // @[PoorAXIL2Reg.scala 31:27]
      s_wr <= 1'h0; // @[PoorAXIL2Reg.scala 31:27]
    end else if (_io_axi_aw_ready_T) begin // @[Conditional.scala 40:58]
      s_wr <= _GEN_1543;
    end else if (s_wr) begin // @[Conditional.scala 39:67]
      if (_T_4) begin // @[PoorAXIL2Reg.scala 75:39]
        s_wr <= 1'h0; // @[PoorAXIL2Reg.scala 76:57]
      end
    end
    if (_io_axi_ar_ready_T) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[PoorAXIL2Reg.scala 50:40]
        r_addr <= _r_addr_T; // @[PoorAXIL2Reg.scala 51:57]
      end
    end
    if (_io_axi_aw_ready_T) begin // @[Conditional.scala 40:58]
      if (_T_7) begin // @[PoorAXIL2Reg.scala 69:40]
        w_addr <= _w_addr_T; // @[PoorAXIL2Reg.scala 70:57]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_control_8 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_control_9 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_control_10 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_control_11 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_control_12 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_control_13 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_control_20 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_control_50 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_control_51 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_control_52 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_control_53 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_control_54 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_control_55 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_control_56 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  reg_control_57 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  reg_control_58 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  reg_control_59 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  reg_control_70 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  reg_control_71 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_control_72 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_control_73 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_control_74 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_control_75 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_control_76 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_control_77 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_control_78 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_control_79 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_control_80 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_control_91 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_control_92 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_control_93 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_control_94 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  reg_status_40 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  reg_status_51 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  reg_status_52 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  reg_status_61 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  reg_status_71 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  reg_status_72 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  reg_status_75 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  reg_status_76 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  reg_status_77 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  reg_status_78 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  reg_status_79 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  reg_status_81 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  s_rd = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  s_wr = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  r_addr = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  w_addr = _RAND_47[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_2(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [511:0] io_enq_bits_data,
  input  [31:0]  io_enq_bits_ctrl_len,
  input          io_enq_bits_last,
  input          io_deq_ready,
  output         io_deq_valid,
  output [511:0] io_deq_bits_data,
  output [31:0]  io_deq_bits_tcrc,
  output         io_deq_bits_ctrl_marker,
  output [6:0]   io_deq_bits_ctrl_ecc,
  output [31:0]  io_deq_bits_ctrl_len,
  output [2:0]   io_deq_bits_ctrl_port_id,
  output [10:0]  io_deq_bits_ctrl_qid,
  output         io_deq_bits_ctrl_has_cmpt,
  output         io_deq_bits_last,
  output [5:0]   io_deq_bits_mty
);
`ifdef RANDOMIZE_MEM_INIT
  reg [511:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] ram_data [0:15]; // @[Decoupled.scala 218:16]
  wire [511:0] ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_data_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [511:0] ram_data_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_data_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_data_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_tcrc [0:15]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_tcrc_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_tcrc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_tcrc_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_tcrc_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_tcrc_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_tcrc_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_ctrl_marker [0:15]; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_marker_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_marker_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_marker_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_marker_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_marker_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_marker_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_ctrl_ecc [0:15]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_ctrl_ecc_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_ecc_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_ctrl_ecc_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_ecc_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_ecc_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_ecc_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_ctrl_len [0:15]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_ctrl_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_ctrl_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_ctrl_port_id [0:15]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_ctrl_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_port_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_ctrl_port_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_port_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_port_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_port_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] ram_ctrl_qid [0:15]; // @[Decoupled.scala 218:16]
  wire [10:0] ram_ctrl_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_qid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [10:0] ram_ctrl_qid_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_qid_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_qid_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_qid_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_ctrl_has_cmpt [0:15]; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_has_cmpt_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_has_cmpt_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_has_cmpt_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_ctrl_has_cmpt_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_has_cmpt_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_ctrl_has_cmpt_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_last [0:15]; // @[Decoupled.scala 218:16]
  wire  ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_last_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_last_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_last_MPORT_en; // @[Decoupled.scala 218:16]
  reg [5:0] ram_mty [0:15]; // @[Decoupled.scala 218:16]
  wire [5:0] ram_mty_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mty_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [5:0] ram_mty_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_mty_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_mty_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_mty_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  assign ram_data_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_data_io_deq_bits_MPORT_data = ram_data[ram_data_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_data_MPORT_data = io_enq_bits_data;
  assign ram_data_MPORT_addr = enq_ptr_value;
  assign ram_data_MPORT_mask = 1'h1;
  assign ram_data_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tcrc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_tcrc_io_deq_bits_MPORT_data = ram_tcrc[ram_tcrc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_tcrc_MPORT_data = 32'h0;
  assign ram_tcrc_MPORT_addr = enq_ptr_value;
  assign ram_tcrc_MPORT_mask = 1'h1;
  assign ram_tcrc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_marker_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_marker_io_deq_bits_MPORT_data = ram_ctrl_marker[ram_ctrl_marker_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_marker_MPORT_data = 1'h0;
  assign ram_ctrl_marker_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_marker_MPORT_mask = 1'h1;
  assign ram_ctrl_marker_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_ecc_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_ecc_io_deq_bits_MPORT_data = ram_ctrl_ecc[ram_ctrl_ecc_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_ecc_MPORT_data = 7'h0;
  assign ram_ctrl_ecc_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_ecc_MPORT_mask = 1'h1;
  assign ram_ctrl_ecc_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_len_io_deq_bits_MPORT_data = ram_ctrl_len[ram_ctrl_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_len_MPORT_data = io_enq_bits_ctrl_len;
  assign ram_ctrl_len_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_len_MPORT_mask = 1'h1;
  assign ram_ctrl_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_port_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_port_id_io_deq_bits_MPORT_data = ram_ctrl_port_id[ram_ctrl_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_port_id_MPORT_data = 3'h0;
  assign ram_ctrl_port_id_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_port_id_MPORT_mask = 1'h1;
  assign ram_ctrl_port_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_qid_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_qid_io_deq_bits_MPORT_data = ram_ctrl_qid[ram_ctrl_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_qid_MPORT_data = 11'h0;
  assign ram_ctrl_qid_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_qid_MPORT_mask = 1'h1;
  assign ram_ctrl_qid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_ctrl_has_cmpt_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_ctrl_has_cmpt_io_deq_bits_MPORT_data = ram_ctrl_has_cmpt[ram_ctrl_has_cmpt_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_ctrl_has_cmpt_MPORT_data = 1'h0;
  assign ram_ctrl_has_cmpt_MPORT_addr = enq_ptr_value;
  assign ram_ctrl_has_cmpt_MPORT_mask = 1'h1;
  assign ram_ctrl_has_cmpt_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_last_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_last_io_deq_bits_MPORT_data = ram_last[ram_last_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_last_MPORT_data = io_enq_bits_last;
  assign ram_last_MPORT_addr = enq_ptr_value;
  assign ram_last_MPORT_mask = 1'h1;
  assign ram_last_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_mty_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_mty_io_deq_bits_MPORT_data = ram_mty[ram_mty_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_mty_MPORT_data = 6'h0;
  assign ram_mty_MPORT_addr = enq_ptr_value;
  assign ram_mty_MPORT_mask = 1'h1;
  assign ram_mty_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_data = ram_data_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_tcrc = ram_tcrc_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_marker = ram_ctrl_marker_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_ecc = ram_ctrl_ecc_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_len = ram_ctrl_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_port_id = ram_ctrl_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_qid = ram_ctrl_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_ctrl_has_cmpt = ram_ctrl_has_cmpt_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_last = ram_last_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_mty = ram_mty_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_data_MPORT_en & ram_data_MPORT_mask) begin
      ram_data[ram_data_MPORT_addr] <= ram_data_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_tcrc_MPORT_en & ram_tcrc_MPORT_mask) begin
      ram_tcrc[ram_tcrc_MPORT_addr] <= ram_tcrc_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_marker_MPORT_en & ram_ctrl_marker_MPORT_mask) begin
      ram_ctrl_marker[ram_ctrl_marker_MPORT_addr] <= ram_ctrl_marker_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_ecc_MPORT_en & ram_ctrl_ecc_MPORT_mask) begin
      ram_ctrl_ecc[ram_ctrl_ecc_MPORT_addr] <= ram_ctrl_ecc_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_len_MPORT_en & ram_ctrl_len_MPORT_mask) begin
      ram_ctrl_len[ram_ctrl_len_MPORT_addr] <= ram_ctrl_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_port_id_MPORT_en & ram_ctrl_port_id_MPORT_mask) begin
      ram_ctrl_port_id[ram_ctrl_port_id_MPORT_addr] <= ram_ctrl_port_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_qid_MPORT_en & ram_ctrl_qid_MPORT_mask) begin
      ram_ctrl_qid[ram_ctrl_qid_MPORT_addr] <= ram_ctrl_qid_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_ctrl_has_cmpt_MPORT_en & ram_ctrl_has_cmpt_MPORT_mask) begin
      ram_ctrl_has_cmpt[ram_ctrl_has_cmpt_MPORT_addr] <= ram_ctrl_has_cmpt_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_last_MPORT_en & ram_last_MPORT_mask) begin
      ram_last[ram_last_MPORT_addr] <= ram_last_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_mty_MPORT_en & ram_mty_MPORT_mask) begin
      ram_mty[ram_mty_MPORT_addr] <= ram_mty_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {16{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_data[initvar] = _RAND_0[511:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_tcrc[initvar] = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_marker[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_ecc[initvar] = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_len[initvar] = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_port_id[initvar] = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_qid[initvar] = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_ctrl_has_cmpt[initvar] = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_last[initvar] = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_mty[initvar] = _RAND_9[5:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  enq_ptr_value = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  deq_ptr_value = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  maybe_full = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [511:0] io_in_bits_data,
  input  [31:0]  io_in_bits_ctrl_len,
  input          io_in_bits_last,
  input          io_out_ready,
  output         io_out_valid,
  output [511:0] io_out_bits_data,
  output [31:0]  io_out_bits_tcrc,
  output         io_out_bits_ctrl_marker,
  output [6:0]   io_out_bits_ctrl_ecc,
  output [31:0]  io_out_bits_ctrl_len,
  output [2:0]   io_out_bits_ctrl_port_id,
  output [10:0]  io_out_bits_ctrl_qid,
  output         io_out_bits_ctrl_has_cmpt,
  output         io_out_bits_last,
  output [5:0]   io_out_bits_mty
);
  wire  q_clock; // @[XQueue.scala 85:39]
  wire  q_reset; // @[XQueue.scala 85:39]
  wire  q_io_enq_ready; // @[XQueue.scala 85:39]
  wire  q_io_enq_valid; // @[XQueue.scala 85:39]
  wire [511:0] q_io_enq_bits_data; // @[XQueue.scala 85:39]
  wire [31:0] q_io_enq_bits_ctrl_len; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_last; // @[XQueue.scala 85:39]
  wire  q_io_deq_ready; // @[XQueue.scala 85:39]
  wire  q_io_deq_valid; // @[XQueue.scala 85:39]
  wire [511:0] q_io_deq_bits_data; // @[XQueue.scala 85:39]
  wire [31:0] q_io_deq_bits_tcrc; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_ctrl_marker; // @[XQueue.scala 85:39]
  wire [6:0] q_io_deq_bits_ctrl_ecc; // @[XQueue.scala 85:39]
  wire [31:0] q_io_deq_bits_ctrl_len; // @[XQueue.scala 85:39]
  wire [2:0] q_io_deq_bits_ctrl_port_id; // @[XQueue.scala 85:39]
  wire [10:0] q_io_deq_bits_ctrl_qid; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_ctrl_has_cmpt; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_last; // @[XQueue.scala 85:39]
  wire [5:0] q_io_deq_bits_mty; // @[XQueue.scala 85:39]
  Queue_2 q ( // @[XQueue.scala 85:39]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_data(q_io_enq_bits_data),
    .io_enq_bits_ctrl_len(q_io_enq_bits_ctrl_len),
    .io_enq_bits_last(q_io_enq_bits_last),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_data(q_io_deq_bits_data),
    .io_deq_bits_tcrc(q_io_deq_bits_tcrc),
    .io_deq_bits_ctrl_marker(q_io_deq_bits_ctrl_marker),
    .io_deq_bits_ctrl_ecc(q_io_deq_bits_ctrl_ecc),
    .io_deq_bits_ctrl_len(q_io_deq_bits_ctrl_len),
    .io_deq_bits_ctrl_port_id(q_io_deq_bits_ctrl_port_id),
    .io_deq_bits_ctrl_qid(q_io_deq_bits_ctrl_qid),
    .io_deq_bits_ctrl_has_cmpt(q_io_deq_bits_ctrl_has_cmpt),
    .io_deq_bits_last(q_io_deq_bits_last),
    .io_deq_bits_mty(q_io_deq_bits_mty)
  );
  assign io_in_ready = q_io_enq_ready; // @[XQueue.scala 87:34]
  assign io_out_valid = q_io_deq_valid; // @[XQueue.scala 88:34]
  assign io_out_bits_data = q_io_deq_bits_data; // @[XQueue.scala 88:34]
  assign io_out_bits_tcrc = q_io_deq_bits_tcrc; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_marker = q_io_deq_bits_ctrl_marker; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_ecc = q_io_deq_bits_ctrl_ecc; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_len = q_io_deq_bits_ctrl_len; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_port_id = q_io_deq_bits_ctrl_port_id; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_qid = q_io_deq_bits_ctrl_qid; // @[XQueue.scala 88:34]
  assign io_out_bits_ctrl_has_cmpt = q_io_deq_bits_ctrl_has_cmpt; // @[XQueue.scala 88:34]
  assign io_out_bits_last = q_io_deq_bits_last; // @[XQueue.scala 88:34]
  assign io_out_bits_mty = q_io_deq_bits_mty; // @[XQueue.scala 88:34]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_valid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_data = io_in_bits_data; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_ctrl_len = io_in_bits_ctrl_len; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_last = io_in_bits_last; // @[XQueue.scala 87:34]
  assign q_io_deq_ready = io_out_ready; // @[XQueue.scala 88:34]
endmodule
module Queue_3(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_addr,
  input  [10:0] io_enq_bits_qid,
  input         io_enq_bits_error,
  input  [7:0]  io_enq_bits_func,
  input  [2:0]  io_enq_bits_port_id,
  input  [6:0]  io_enq_bits_pfch_tag,
  input  [31:0] io_enq_bits_len,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_addr,
  output [10:0] io_deq_bits_qid,
  output        io_deq_bits_error,
  output [7:0]  io_deq_bits_func,
  output [2:0]  io_deq_bits_port_id,
  output [6:0]  io_deq_bits_pfch_tag,
  output [31:0] io_deq_bits_len
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_addr [0:15]; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [63:0] ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_addr_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 218:16]
  reg [10:0] ram_qid [0:15]; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [10:0] ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_qid_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_qid_MPORT_en; // @[Decoupled.scala 218:16]
  reg  ram_error [0:15]; // @[Decoupled.scala 218:16]
  wire  ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_error_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_error_MPORT_en; // @[Decoupled.scala 218:16]
  reg [7:0] ram_func [0:15]; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [7:0] ram_func_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_func_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_func_MPORT_en; // @[Decoupled.scala 218:16]
  reg [2:0] ram_port_id [0:15]; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [2:0] ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_port_id_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_port_id_MPORT_en; // @[Decoupled.scala 218:16]
  reg [6:0] ram_pfch_tag [0:15]; // @[Decoupled.scala 218:16]
  wire [6:0] ram_pfch_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_pfch_tag_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [6:0] ram_pfch_tag_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_pfch_tag_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_pfch_tag_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_pfch_tag_MPORT_en; // @[Decoupled.scala 218:16]
  reg [31:0] ram_len [0:15]; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [31:0] ram_len_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_len_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  assign ram_addr_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = enq_ptr_value;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_qid_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_qid_io_deq_bits_MPORT_data = ram_qid[ram_qid_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_qid_MPORT_data = io_enq_bits_qid;
  assign ram_qid_MPORT_addr = enq_ptr_value;
  assign ram_qid_MPORT_mask = 1'h1;
  assign ram_qid_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_error_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_error_io_deq_bits_MPORT_data = ram_error[ram_error_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_error_MPORT_data = io_enq_bits_error;
  assign ram_error_MPORT_addr = enq_ptr_value;
  assign ram_error_MPORT_mask = 1'h1;
  assign ram_error_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_func_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_func_io_deq_bits_MPORT_data = ram_func[ram_func_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_func_MPORT_data = io_enq_bits_func;
  assign ram_func_MPORT_addr = enq_ptr_value;
  assign ram_func_MPORT_mask = 1'h1;
  assign ram_func_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_port_id_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_port_id_io_deq_bits_MPORT_data = ram_port_id[ram_port_id_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_port_id_MPORT_data = io_enq_bits_port_id;
  assign ram_port_id_MPORT_addr = enq_ptr_value;
  assign ram_port_id_MPORT_mask = 1'h1;
  assign ram_port_id_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_pfch_tag_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_pfch_tag_io_deq_bits_MPORT_data = ram_pfch_tag[ram_pfch_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_pfch_tag_MPORT_data = io_enq_bits_pfch_tag;
  assign ram_pfch_tag_MPORT_addr = enq_ptr_value;
  assign ram_pfch_tag_MPORT_mask = 1'h1;
  assign ram_pfch_tag_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = enq_ptr_value;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_qid = ram_qid_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_error = ram_error_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_func = ram_func_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_port_id = ram_port_id_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_pfch_tag = ram_pfch_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_qid_MPORT_en & ram_qid_MPORT_mask) begin
      ram_qid[ram_qid_MPORT_addr] <= ram_qid_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_error_MPORT_en & ram_error_MPORT_mask) begin
      ram_error[ram_error_MPORT_addr] <= ram_error_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_func_MPORT_en & ram_func_MPORT_mask) begin
      ram_func[ram_func_MPORT_addr] <= ram_func_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_port_id_MPORT_en & ram_port_id_MPORT_mask) begin
      ram_port_id[ram_port_id_MPORT_addr] <= ram_port_id_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_pfch_tag_MPORT_en & ram_pfch_tag_MPORT_mask) begin
      ram_pfch_tag[ram_pfch_tag_MPORT_addr] <= ram_pfch_tag_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if(ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_qid[initvar] = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_error[initvar] = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_func[initvar] = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_port_id[initvar] = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_pfch_tag[initvar] = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_len[initvar] = _RAND_6[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  enq_ptr_value = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  deq_ptr_value = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  maybe_full = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_addr,
  input  [10:0] io_in_bits_qid,
  input         io_in_bits_error,
  input  [7:0]  io_in_bits_func,
  input  [2:0]  io_in_bits_port_id,
  input  [6:0]  io_in_bits_pfch_tag,
  input  [31:0] io_in_bits_len,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_addr,
  output [10:0] io_out_bits_qid,
  output        io_out_bits_error,
  output [7:0]  io_out_bits_func,
  output [2:0]  io_out_bits_port_id,
  output [6:0]  io_out_bits_pfch_tag,
  output [31:0] io_out_bits_len
);
  wire  q_clock; // @[XQueue.scala 85:39]
  wire  q_reset; // @[XQueue.scala 85:39]
  wire  q_io_enq_ready; // @[XQueue.scala 85:39]
  wire  q_io_enq_valid; // @[XQueue.scala 85:39]
  wire [63:0] q_io_enq_bits_addr; // @[XQueue.scala 85:39]
  wire [10:0] q_io_enq_bits_qid; // @[XQueue.scala 85:39]
  wire  q_io_enq_bits_error; // @[XQueue.scala 85:39]
  wire [7:0] q_io_enq_bits_func; // @[XQueue.scala 85:39]
  wire [2:0] q_io_enq_bits_port_id; // @[XQueue.scala 85:39]
  wire [6:0] q_io_enq_bits_pfch_tag; // @[XQueue.scala 85:39]
  wire [31:0] q_io_enq_bits_len; // @[XQueue.scala 85:39]
  wire  q_io_deq_ready; // @[XQueue.scala 85:39]
  wire  q_io_deq_valid; // @[XQueue.scala 85:39]
  wire [63:0] q_io_deq_bits_addr; // @[XQueue.scala 85:39]
  wire [10:0] q_io_deq_bits_qid; // @[XQueue.scala 85:39]
  wire  q_io_deq_bits_error; // @[XQueue.scala 85:39]
  wire [7:0] q_io_deq_bits_func; // @[XQueue.scala 85:39]
  wire [2:0] q_io_deq_bits_port_id; // @[XQueue.scala 85:39]
  wire [6:0] q_io_deq_bits_pfch_tag; // @[XQueue.scala 85:39]
  wire [31:0] q_io_deq_bits_len; // @[XQueue.scala 85:39]
  Queue_3 q ( // @[XQueue.scala 85:39]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits_addr(q_io_enq_bits_addr),
    .io_enq_bits_qid(q_io_enq_bits_qid),
    .io_enq_bits_error(q_io_enq_bits_error),
    .io_enq_bits_func(q_io_enq_bits_func),
    .io_enq_bits_port_id(q_io_enq_bits_port_id),
    .io_enq_bits_pfch_tag(q_io_enq_bits_pfch_tag),
    .io_enq_bits_len(q_io_enq_bits_len),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits_addr(q_io_deq_bits_addr),
    .io_deq_bits_qid(q_io_deq_bits_qid),
    .io_deq_bits_error(q_io_deq_bits_error),
    .io_deq_bits_func(q_io_deq_bits_func),
    .io_deq_bits_port_id(q_io_deq_bits_port_id),
    .io_deq_bits_pfch_tag(q_io_deq_bits_pfch_tag),
    .io_deq_bits_len(q_io_deq_bits_len)
  );
  assign io_in_ready = q_io_enq_ready; // @[XQueue.scala 87:34]
  assign io_out_valid = q_io_deq_valid; // @[XQueue.scala 88:34]
  assign io_out_bits_addr = q_io_deq_bits_addr; // @[XQueue.scala 88:34]
  assign io_out_bits_qid = q_io_deq_bits_qid; // @[XQueue.scala 88:34]
  assign io_out_bits_error = q_io_deq_bits_error; // @[XQueue.scala 88:34]
  assign io_out_bits_func = q_io_deq_bits_func; // @[XQueue.scala 88:34]
  assign io_out_bits_port_id = q_io_deq_bits_port_id; // @[XQueue.scala 88:34]
  assign io_out_bits_pfch_tag = q_io_deq_bits_pfch_tag; // @[XQueue.scala 88:34]
  assign io_out_bits_len = q_io_deq_bits_len; // @[XQueue.scala 88:34]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_valid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_addr = io_in_bits_addr; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_qid = io_in_bits_qid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_error = io_in_bits_error; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_func = io_in_bits_func; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_port_id = io_in_bits_port_id; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_pfch_tag = io_in_bits_pfch_tag; // @[XQueue.scala 87:34]
  assign q_io_enq_bits_len = io_in_bits_len; // @[XQueue.scala 87:34]
  assign q_io_deq_ready = io_out_ready; // @[XQueue.scala 88:34]
endmodule
module DataBoundarySplit(
  input          clock,
  input          reset,
  output         io_data_in_ready,
  input          io_data_in_valid,
  input  [511:0] io_data_in_bits_data,
  output         io_cmd_in_ready,
  input          io_cmd_in_valid,
  input  [63:0]  io_cmd_in_bits_addr,
  input  [10:0]  io_cmd_in_bits_qid,
  input          io_cmd_in_bits_error,
  input  [7:0]   io_cmd_in_bits_func,
  input  [2:0]   io_cmd_in_bits_port_id,
  input  [6:0]   io_cmd_in_bits_pfch_tag,
  input  [31:0]  io_cmd_in_bits_len,
  input          io_data_out_ready,
  output         io_data_out_valid,
  output [511:0] io_data_out_bits_data,
  output [31:0]  io_data_out_bits_tcrc,
  output         io_data_out_bits_ctrl_marker,
  output [6:0]   io_data_out_bits_ctrl_ecc,
  output [31:0]  io_data_out_bits_ctrl_len,
  output [2:0]   io_data_out_bits_ctrl_port_id,
  output [10:0]  io_data_out_bits_ctrl_qid,
  output         io_data_out_bits_ctrl_has_cmpt,
  output         io_data_out_bits_last,
  output [5:0]   io_data_out_bits_mty,
  input          io_cmd_out_ready,
  output         io_cmd_out_valid,
  output [63:0]  io_cmd_out_bits_addr,
  output [10:0]  io_cmd_out_bits_qid,
  output         io_cmd_out_bits_error,
  output [7:0]   io_cmd_out_bits_func,
  output [2:0]   io_cmd_out_bits_port_id,
  output [6:0]   io_cmd_out_bits_pfch_tag,
  output [31:0]  io_cmd_out_bits_len
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  data_fifo_clock; // @[XQueue.scala 35:23]
  wire  data_fifo_reset; // @[XQueue.scala 35:23]
  wire  data_fifo_io_in_ready; // @[XQueue.scala 35:23]
  wire  data_fifo_io_in_valid; // @[XQueue.scala 35:23]
  wire [511:0] data_fifo_io_in_bits_data; // @[XQueue.scala 35:23]
  wire [31:0] data_fifo_io_in_bits_ctrl_len; // @[XQueue.scala 35:23]
  wire  data_fifo_io_in_bits_last; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_ready; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_valid; // @[XQueue.scala 35:23]
  wire [511:0] data_fifo_io_out_bits_data; // @[XQueue.scala 35:23]
  wire [31:0] data_fifo_io_out_bits_tcrc; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_bits_ctrl_marker; // @[XQueue.scala 35:23]
  wire [6:0] data_fifo_io_out_bits_ctrl_ecc; // @[XQueue.scala 35:23]
  wire [31:0] data_fifo_io_out_bits_ctrl_len; // @[XQueue.scala 35:23]
  wire [2:0] data_fifo_io_out_bits_ctrl_port_id; // @[XQueue.scala 35:23]
  wire [10:0] data_fifo_io_out_bits_ctrl_qid; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_bits_ctrl_has_cmpt; // @[XQueue.scala 35:23]
  wire  data_fifo_io_out_bits_last; // @[XQueue.scala 35:23]
  wire [5:0] data_fifo_io_out_bits_mty; // @[XQueue.scala 35:23]
  wire  cmd_fifo_clock; // @[XQueue.scala 35:23]
  wire  cmd_fifo_reset; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_in_ready; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] cmd_fifo_io_in_bits_addr; // @[XQueue.scala 35:23]
  wire [10:0] cmd_fifo_io_in_bits_qid; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_in_bits_error; // @[XQueue.scala 35:23]
  wire [7:0] cmd_fifo_io_in_bits_func; // @[XQueue.scala 35:23]
  wire [2:0] cmd_fifo_io_in_bits_port_id; // @[XQueue.scala 35:23]
  wire [6:0] cmd_fifo_io_in_bits_pfch_tag; // @[XQueue.scala 35:23]
  wire [31:0] cmd_fifo_io_in_bits_len; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_out_ready; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] cmd_fifo_io_out_bits_addr; // @[XQueue.scala 35:23]
  wire [10:0] cmd_fifo_io_out_bits_qid; // @[XQueue.scala 35:23]
  wire  cmd_fifo_io_out_bits_error; // @[XQueue.scala 35:23]
  wire [7:0] cmd_fifo_io_out_bits_func; // @[XQueue.scala 35:23]
  wire [2:0] cmd_fifo_io_out_bits_port_id; // @[XQueue.scala 35:23]
  wire [6:0] cmd_fifo_io_out_bits_pfch_tag; // @[XQueue.scala 35:23]
  wire [31:0] cmd_fifo_io_out_bits_len; // @[XQueue.scala 35:23]
  reg [31:0] cmd_temp_len; // @[CheckSplit.scala 22:27]
  reg [31:0] clength; // @[CheckSplit.scala 23:30]
  reg  state; // @[CheckSplit.scala 28:50]
  reg  tmp_reg; // @[CheckSplit.scala 29:42]
  wire  _io_cmd_in_ready_T = ~state; // @[CheckSplit.scala 34:67]
  wire  _T_2 = io_cmd_in_ready & io_cmd_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_8 = _T_2 | state; // @[CheckSplit.scala 47:47 CheckSplit.scala 49:41 CheckSplit.scala 28:50]
  wire [31:0] _GEN_10 = _T_2 ? io_cmd_in_bits_len : 32'h0; // @[CheckSplit.scala 47:47 CheckSplit.scala 51:57 CheckSplit.scala 40:65]
  wire [6:0] _GEN_11 = _T_2 ? io_cmd_in_bits_pfch_tag : 7'h0; // @[CheckSplit.scala 47:47 CheckSplit.scala 51:57 CheckSplit.scala 40:65]
  wire [2:0] _GEN_12 = _T_2 ? io_cmd_in_bits_port_id : 3'h0; // @[CheckSplit.scala 47:47 CheckSplit.scala 51:57 CheckSplit.scala 40:65]
  wire [7:0] _GEN_13 = _T_2 ? io_cmd_in_bits_func : 8'h0; // @[CheckSplit.scala 47:47 CheckSplit.scala 51:57 CheckSplit.scala 40:65]
  wire  _GEN_14 = _T_2 & io_cmd_in_bits_error; // @[CheckSplit.scala 47:47 CheckSplit.scala 51:57 CheckSplit.scala 40:65]
  wire [10:0] _GEN_15 = _T_2 ? io_cmd_in_bits_qid : 11'h0; // @[CheckSplit.scala 47:47 CheckSplit.scala 51:57 CheckSplit.scala 40:65]
  wire [63:0] _GEN_16 = _T_2 ? io_cmd_in_bits_addr : 64'h0; // @[CheckSplit.scala 47:47 CheckSplit.scala 51:57 CheckSplit.scala 40:65]
  wire  _GEN_17 = _T_2 | tmp_reg; // @[CheckSplit.scala 47:47 CheckSplit.scala 52:73 CheckSplit.scala 29:42]
  wire  _T_3 = io_data_in_ready & io_data_in_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _clength_T_1 = clength + 32'h40; // @[CheckSplit.scala 60:100]
  wire  _T_6 = _clength_T_1 >= io_cmd_in_bits_len; // @[CheckSplit.scala 61:55]
  wire  _GEN_25 = _T_3 & _T_6; // @[CheckSplit.scala 55:48 CheckSplit.scala 38:57]
  wire [31:0] _GEN_29 = _T_3 ? io_cmd_in_bits_len : 32'h0; // @[CheckSplit.scala 55:48 CheckSplit.scala 59:65 CheckSplit.scala 38:57]
  wire [511:0] _GEN_33 = _T_3 ? io_data_in_bits_data : 512'h0; // @[CheckSplit.scala 55:48 CheckSplit.scala 57:73 CheckSplit.scala 38:57]
  wire  _T_11 = _clength_T_1 >= cmd_temp_len; // @[CheckSplit.scala 76:55]
  wire  _GEN_38 = _clength_T_1 >= cmd_temp_len ? 1'h0 : state; // @[CheckSplit.scala 76:71 CheckSplit.scala 78:89 CheckSplit.scala 28:50]
  wire  _GEN_39 = _clength_T_1 >= cmd_temp_len ? 1'h0 : tmp_reg; // @[CheckSplit.scala 76:71 CheckSplit.scala 79:89 CheckSplit.scala 29:42]
  wire [31:0] _GEN_40 = _clength_T_1 >= cmd_temp_len ? 32'h0 : _clength_T_1; // @[CheckSplit.scala 76:71 CheckSplit.scala 80:89 CheckSplit.scala 75:89]
  wire  _GEN_43 = _T_3 & _T_11; // @[CheckSplit.scala 70:48 CheckSplit.scala 38:57]
  wire [31:0] _GEN_47 = _T_3 ? cmd_temp_len : 32'h0; // @[CheckSplit.scala 70:48 CheckSplit.scala 74:65 CheckSplit.scala 38:57]
  wire  _GEN_55 = state & _T_3; // @[Conditional.scala 39:67 CheckSplit.scala 37:57]
  wire  _GEN_57 = state & _GEN_43; // @[Conditional.scala 39:67 CheckSplit.scala 38:57]
  wire [31:0] _GEN_61 = state ? _GEN_47 : 32'h0; // @[Conditional.scala 39:67 CheckSplit.scala 38:57]
  wire [511:0] _GEN_65 = state ? _GEN_33 : 512'h0; // @[Conditional.scala 39:67 CheckSplit.scala 38:57]
  XQueue data_fifo ( // @[XQueue.scala 35:23]
    .clock(data_fifo_clock),
    .reset(data_fifo_reset),
    .io_in_ready(data_fifo_io_in_ready),
    .io_in_valid(data_fifo_io_in_valid),
    .io_in_bits_data(data_fifo_io_in_bits_data),
    .io_in_bits_ctrl_len(data_fifo_io_in_bits_ctrl_len),
    .io_in_bits_last(data_fifo_io_in_bits_last),
    .io_out_ready(data_fifo_io_out_ready),
    .io_out_valid(data_fifo_io_out_valid),
    .io_out_bits_data(data_fifo_io_out_bits_data),
    .io_out_bits_tcrc(data_fifo_io_out_bits_tcrc),
    .io_out_bits_ctrl_marker(data_fifo_io_out_bits_ctrl_marker),
    .io_out_bits_ctrl_ecc(data_fifo_io_out_bits_ctrl_ecc),
    .io_out_bits_ctrl_len(data_fifo_io_out_bits_ctrl_len),
    .io_out_bits_ctrl_port_id(data_fifo_io_out_bits_ctrl_port_id),
    .io_out_bits_ctrl_qid(data_fifo_io_out_bits_ctrl_qid),
    .io_out_bits_ctrl_has_cmpt(data_fifo_io_out_bits_ctrl_has_cmpt),
    .io_out_bits_last(data_fifo_io_out_bits_last),
    .io_out_bits_mty(data_fifo_io_out_bits_mty)
  );
  XQueue_1 cmd_fifo ( // @[XQueue.scala 35:23]
    .clock(cmd_fifo_clock),
    .reset(cmd_fifo_reset),
    .io_in_ready(cmd_fifo_io_in_ready),
    .io_in_valid(cmd_fifo_io_in_valid),
    .io_in_bits_addr(cmd_fifo_io_in_bits_addr),
    .io_in_bits_qid(cmd_fifo_io_in_bits_qid),
    .io_in_bits_error(cmd_fifo_io_in_bits_error),
    .io_in_bits_func(cmd_fifo_io_in_bits_func),
    .io_in_bits_port_id(cmd_fifo_io_in_bits_port_id),
    .io_in_bits_pfch_tag(cmd_fifo_io_in_bits_pfch_tag),
    .io_in_bits_len(cmd_fifo_io_in_bits_len),
    .io_out_ready(cmd_fifo_io_out_ready),
    .io_out_valid(cmd_fifo_io_out_valid),
    .io_out_bits_addr(cmd_fifo_io_out_bits_addr),
    .io_out_bits_qid(cmd_fifo_io_out_bits_qid),
    .io_out_bits_error(cmd_fifo_io_out_bits_error),
    .io_out_bits_func(cmd_fifo_io_out_bits_func),
    .io_out_bits_port_id(cmd_fifo_io_out_bits_port_id),
    .io_out_bits_pfch_tag(cmd_fifo_io_out_bits_pfch_tag),
    .io_out_bits_len(cmd_fifo_io_out_bits_len)
  );
  assign io_data_in_ready = data_fifo_io_in_ready & tmp_reg; // @[CheckSplit.scala 35:92]
  assign io_cmd_in_ready = ~state & cmd_fifo_io_in_ready; // @[CheckSplit.scala 34:78]
  assign io_data_out_valid = data_fifo_io_out_valid; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_data = data_fifo_io_out_bits_data; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_tcrc = data_fifo_io_out_bits_tcrc; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_ctrl_marker = data_fifo_io_out_bits_ctrl_marker; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_ctrl_ecc = data_fifo_io_out_bits_ctrl_ecc; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_ctrl_len = data_fifo_io_out_bits_ctrl_len; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_ctrl_port_id = data_fifo_io_out_bits_ctrl_port_id; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_ctrl_qid = data_fifo_io_out_bits_ctrl_qid; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_ctrl_has_cmpt = data_fifo_io_out_bits_ctrl_has_cmpt; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_last = data_fifo_io_out_bits_last; // @[CheckSplit.scala 24:25]
  assign io_data_out_bits_mty = data_fifo_io_out_bits_mty; // @[CheckSplit.scala 24:25]
  assign io_cmd_out_valid = cmd_fifo_io_out_valid; // @[CheckSplit.scala 25:25]
  assign io_cmd_out_bits_addr = cmd_fifo_io_out_bits_addr; // @[CheckSplit.scala 25:25]
  assign io_cmd_out_bits_qid = cmd_fifo_io_out_bits_qid; // @[CheckSplit.scala 25:25]
  assign io_cmd_out_bits_error = cmd_fifo_io_out_bits_error; // @[CheckSplit.scala 25:25]
  assign io_cmd_out_bits_func = cmd_fifo_io_out_bits_func; // @[CheckSplit.scala 25:25]
  assign io_cmd_out_bits_port_id = cmd_fifo_io_out_bits_port_id; // @[CheckSplit.scala 25:25]
  assign io_cmd_out_bits_pfch_tag = cmd_fifo_io_out_bits_pfch_tag; // @[CheckSplit.scala 25:25]
  assign io_cmd_out_bits_len = cmd_fifo_io_out_bits_len; // @[CheckSplit.scala 25:25]
  assign data_fifo_clock = clock;
  assign data_fifo_reset = reset;
  assign data_fifo_io_in_valid = _io_cmd_in_ready_T ? _T_3 : _GEN_55; // @[Conditional.scala 40:58]
  assign data_fifo_io_in_bits_data = _io_cmd_in_ready_T ? _GEN_33 : _GEN_65; // @[Conditional.scala 40:58]
  assign data_fifo_io_in_bits_ctrl_len = _io_cmd_in_ready_T ? _GEN_29 : _GEN_61; // @[Conditional.scala 40:58]
  assign data_fifo_io_in_bits_last = _io_cmd_in_ready_T ? _GEN_25 : _GEN_57; // @[Conditional.scala 40:58]
  assign data_fifo_io_out_ready = io_data_out_ready; // @[CheckSplit.scala 24:25]
  assign cmd_fifo_clock = clock;
  assign cmd_fifo_reset = reset;
  assign cmd_fifo_io_in_valid = _io_cmd_in_ready_T & _T_2; // @[Conditional.scala 40:58 CheckSplit.scala 39:57]
  assign cmd_fifo_io_in_bits_addr = _io_cmd_in_ready_T ? _GEN_16 : 64'h0; // @[Conditional.scala 40:58 CheckSplit.scala 40:65]
  assign cmd_fifo_io_in_bits_qid = _io_cmd_in_ready_T ? _GEN_15 : 11'h0; // @[Conditional.scala 40:58 CheckSplit.scala 40:65]
  assign cmd_fifo_io_in_bits_error = _io_cmd_in_ready_T & _GEN_14; // @[Conditional.scala 40:58 CheckSplit.scala 40:65]
  assign cmd_fifo_io_in_bits_func = _io_cmd_in_ready_T ? _GEN_13 : 8'h0; // @[Conditional.scala 40:58 CheckSplit.scala 40:65]
  assign cmd_fifo_io_in_bits_port_id = _io_cmd_in_ready_T ? _GEN_12 : 3'h0; // @[Conditional.scala 40:58 CheckSplit.scala 40:65]
  assign cmd_fifo_io_in_bits_pfch_tag = _io_cmd_in_ready_T ? _GEN_11 : 7'h0; // @[Conditional.scala 40:58 CheckSplit.scala 40:65]
  assign cmd_fifo_io_in_bits_len = _io_cmd_in_ready_T ? _GEN_10 : 32'h0; // @[Conditional.scala 40:58 CheckSplit.scala 40:65]
  assign cmd_fifo_io_out_ready = io_cmd_out_ready; // @[CheckSplit.scala 25:25]
  always @(posedge clock) begin
    if (_io_cmd_in_ready_T) begin // @[Conditional.scala 40:58]
      if (_T_2) begin // @[CheckSplit.scala 47:47]
        cmd_temp_len <= io_cmd_in_bits_len; // @[CheckSplit.scala 48:73]
      end
    end
    if (reset) begin // @[CheckSplit.scala 23:30]
      clength <= 32'h0; // @[CheckSplit.scala 23:30]
    end else if (_io_cmd_in_ready_T) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[CheckSplit.scala 55:48]
        if (_clength_T_1 >= io_cmd_in_bits_len) begin // @[CheckSplit.scala 61:77]
          clength <= 32'h0; // @[CheckSplit.scala 65:89]
        end else begin
          clength <= _clength_T_1; // @[CheckSplit.scala 60:89]
        end
      end
    end else if (state) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[CheckSplit.scala 70:48]
        clength <= _GEN_40;
      end
    end
    if (reset) begin // @[CheckSplit.scala 28:50]
      state <= 1'h0; // @[CheckSplit.scala 28:50]
    end else if (_io_cmd_in_ready_T) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[CheckSplit.scala 55:48]
        if (_clength_T_1 >= io_cmd_in_bits_len) begin // @[CheckSplit.scala 61:77]
          state <= 1'h0; // @[CheckSplit.scala 63:89]
        end else begin
          state <= _GEN_8;
        end
      end else begin
        state <= _GEN_8;
      end
    end else if (state) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[CheckSplit.scala 70:48]
        state <= _GEN_38;
      end
    end
    if (reset) begin // @[CheckSplit.scala 29:42]
      tmp_reg <= 1'h0; // @[CheckSplit.scala 29:42]
    end else if (_io_cmd_in_ready_T) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[CheckSplit.scala 55:48]
        if (_clength_T_1 >= io_cmd_in_bits_len) begin // @[CheckSplit.scala 61:77]
          tmp_reg <= 1'h0; // @[CheckSplit.scala 64:89]
        end else begin
          tmp_reg <= _GEN_17;
        end
      end else begin
        tmp_reg <= _GEN_17;
      end
    end else if (state) begin // @[Conditional.scala 39:67]
      if (_T_3) begin // @[CheckSplit.scala 70:48]
        tmp_reg <= _GEN_39;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmd_temp_len = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  clength = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  tmp_reg = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module QDMA(
  output [15:0]  io_pin_tx_p,
  output [15:0]  io_pin_tx_n,
  input  [15:0]  io_pin_rx_p,
  input  [15:0]  io_pin_rx_n,
  input          io_pin_sys_clk_p,
  input          io_pin_sys_clk_n,
  input          io_pin_sys_rst_n,
  output         io_pcie_clk,
  output         io_pcie_arstn,
  input          io_user_clk,
  input          io_user_arstn,
  output         io_h2c_cmd_ready,
  input          io_h2c_cmd_valid,
  input  [63:0]  io_h2c_cmd_bits_addr,
  input  [31:0]  io_h2c_cmd_bits_len,
  input          io_h2c_data_ready,
  output         io_h2c_data_valid,
  output [511:0] io_h2c_data_bits_data,
  output         io_c2h_cmd_ready,
  input          io_c2h_cmd_valid,
  input  [63:0]  io_c2h_cmd_bits_addr,
  input  [6:0]   io_c2h_cmd_bits_pfch_tag,
  input  [31:0]  io_c2h_cmd_bits_len,
  output         io_c2h_data_ready,
  input          io_c2h_data_valid,
  input  [511:0] io_c2h_data_bits_data,
  output [31:0]  io_reg_control_8,
  output [31:0]  io_reg_control_9,
  output [31:0]  io_reg_control_10,
  output [31:0]  io_reg_control_11,
  output [31:0]  io_reg_control_12,
  output [31:0]  io_reg_control_13,
  output [31:0]  io_reg_control_20,
  output [31:0]  io_reg_control_50,
  output [31:0]  io_reg_control_51,
  output [31:0]  io_reg_control_52,
  output [31:0]  io_reg_control_53,
  output [31:0]  io_reg_control_54,
  output [31:0]  io_reg_control_55,
  output [31:0]  io_reg_control_56,
  output [31:0]  io_reg_control_57,
  output [31:0]  io_reg_control_58,
  output [31:0]  io_reg_control_59,
  output [31:0]  io_reg_control_70,
  output [31:0]  io_reg_control_71,
  output [31:0]  io_reg_control_72,
  output [31:0]  io_reg_control_73,
  output [31:0]  io_reg_control_74,
  output [31:0]  io_reg_control_75,
  output [31:0]  io_reg_control_76,
  output [31:0]  io_reg_control_77,
  output [31:0]  io_reg_control_78,
  output [31:0]  io_reg_control_79,
  output [31:0]  io_reg_control_80,
  output [31:0]  io_reg_control_91,
  output [31:0]  io_reg_control_92,
  output [31:0]  io_reg_control_93,
  output [31:0]  io_reg_control_94,
  input  [31:0]  io_reg_status_40,
  input  [31:0]  io_reg_status_51,
  input  [31:0]  io_reg_status_52,
  input  [31:0]  io_reg_status_61,
  input  [31:0]  io_reg_status_71,
  input  [31:0]  io_reg_status_72,
  input  [31:0]  io_reg_status_75,
  input  [31:0]  io_reg_status_76,
  input  [31:0]  io_reg_status_77,
  input  [31:0]  io_reg_status_78,
  input  [31:0]  io_reg_status_79,
  input  [31:0]  io_reg_status_81,
  input          io_axib_aw_ready,
  output         io_axib_aw_valid,
  output [63:0]  io_axib_aw_bits_addr,
  output [1:0]   io_axib_aw_bits_burst,
  output [7:0]   io_axib_aw_bits_len,
  output [2:0]   io_axib_aw_bits_size,
  input          io_axib_ar_ready,
  output         io_axib_ar_valid,
  output [63:0]  io_axib_ar_bits_addr,
  output [1:0]   io_axib_ar_bits_burst,
  output [7:0]   io_axib_ar_bits_len,
  output [2:0]   io_axib_ar_bits_size,
  input          io_axib_w_ready,
  output         io_axib_w_valid,
  output [511:0] io_axib_w_bits_data,
  output         io_axib_w_bits_last,
  output [63:0]  io_axib_w_bits_strb,
  output         io_axib_r_ready,
  input          io_axib_r_valid,
  input  [511:0] io_axib_r_bits_data,
  input          io_axib_r_bits_last,
  input          io_axib_b_valid,
  output         io_c2h_status_last,
  output         io_c2h_status_cmp,
  output         io_c2h_status_valid,
  output         io_c2h_status_error,
  output         io_c2h_status_drop,
  output [31:0]  io_tlb_miss_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  perst_n_pad_O; // @[Buf.scala 17:34]
  wire  perst_n_pad_I; // @[Buf.scala 17:34]
  wire  ibufds_gte4_inst_O; // @[QDMA.scala 70:38]
  wire  ibufds_gte4_inst_ODIV2; // @[QDMA.scala 70:38]
  wire  ibufds_gte4_inst_CEB; // @[QDMA.scala 70:38]
  wire  ibufds_gte4_inst_I; // @[QDMA.scala 70:38]
  wire  ibufds_gte4_inst_IB; // @[QDMA.scala 70:38]
  wire  fifo_h2c_data_io_in_clk; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_out_clk; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_rstn; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_in_ready; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_in_valid; // @[XConverter.scala 61:33]
  wire [511:0] fifo_h2c_data_io_in_bits_data; // @[XConverter.scala 61:33]
  wire [31:0] fifo_h2c_data_io_in_bits_tcrc; // @[XConverter.scala 61:33]
  wire [10:0] fifo_h2c_data_io_in_bits_tuser_qid; // @[XConverter.scala 61:33]
  wire [2:0] fifo_h2c_data_io_in_bits_tuser_port_id; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_in_bits_tuser_err; // @[XConverter.scala 61:33]
  wire [31:0] fifo_h2c_data_io_in_bits_tuser_mdata; // @[XConverter.scala 61:33]
  wire [5:0] fifo_h2c_data_io_in_bits_tuser_mty; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_in_bits_tuser_zero_byte; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_in_bits_last; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_out_ready; // @[XConverter.scala 61:33]
  wire  fifo_h2c_data_io_out_valid; // @[XConverter.scala 61:33]
  wire [511:0] fifo_h2c_data_io_out_bits_data; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_in_clk; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_out_clk; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_rstn; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_in_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_in_valid; // @[XConverter.scala 61:33]
  wire [511:0] fifo_c2h_data_io_in_bits_data; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_data_io_in_bits_tcrc; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_in_bits_ctrl_marker; // @[XConverter.scala 61:33]
  wire [6:0] fifo_c2h_data_io_in_bits_ctrl_ecc; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_data_io_in_bits_ctrl_len; // @[XConverter.scala 61:33]
  wire [2:0] fifo_c2h_data_io_in_bits_ctrl_port_id; // @[XConverter.scala 61:33]
  wire [10:0] fifo_c2h_data_io_in_bits_ctrl_qid; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_in_bits_ctrl_has_cmpt; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_in_bits_last; // @[XConverter.scala 61:33]
  wire [5:0] fifo_c2h_data_io_in_bits_mty; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_out_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_out_valid; // @[XConverter.scala 61:33]
  wire [511:0] fifo_c2h_data_io_out_bits_data; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_data_io_out_bits_tcrc; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_out_bits_ctrl_marker; // @[XConverter.scala 61:33]
  wire [6:0] fifo_c2h_data_io_out_bits_ctrl_ecc; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_data_io_out_bits_ctrl_len; // @[XConverter.scala 61:33]
  wire [2:0] fifo_c2h_data_io_out_bits_ctrl_port_id; // @[XConverter.scala 61:33]
  wire [10:0] fifo_c2h_data_io_out_bits_ctrl_qid; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_out_bits_ctrl_has_cmpt; // @[XConverter.scala 61:33]
  wire  fifo_c2h_data_io_out_bits_last; // @[XConverter.scala 61:33]
  wire [5:0] fifo_c2h_data_io_out_bits_mty; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_clk; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_clk; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_rstn; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_ready; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_valid; // @[XConverter.scala 61:33]
  wire [63:0] fifo_h2c_cmd_io_in_bits_addr; // @[XConverter.scala 61:33]
  wire [31:0] fifo_h2c_cmd_io_in_bits_len; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_bits_eop; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_bits_sop; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_bits_mrkr_req; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_bits_sdi; // @[XConverter.scala 61:33]
  wire [10:0] fifo_h2c_cmd_io_in_bits_qid; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_bits_error; // @[XConverter.scala 61:33]
  wire [7:0] fifo_h2c_cmd_io_in_bits_func; // @[XConverter.scala 61:33]
  wire [15:0] fifo_h2c_cmd_io_in_bits_cidx; // @[XConverter.scala 61:33]
  wire [2:0] fifo_h2c_cmd_io_in_bits_port_id; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_in_bits_no_dma; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_ready; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_valid; // @[XConverter.scala 61:33]
  wire [63:0] fifo_h2c_cmd_io_out_bits_addr; // @[XConverter.scala 61:33]
  wire [31:0] fifo_h2c_cmd_io_out_bits_len; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_bits_eop; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_bits_sop; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_bits_mrkr_req; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_bits_sdi; // @[XConverter.scala 61:33]
  wire [10:0] fifo_h2c_cmd_io_out_bits_qid; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_bits_error; // @[XConverter.scala 61:33]
  wire [7:0] fifo_h2c_cmd_io_out_bits_func; // @[XConverter.scala 61:33]
  wire [15:0] fifo_h2c_cmd_io_out_bits_cidx; // @[XConverter.scala 61:33]
  wire [2:0] fifo_h2c_cmd_io_out_bits_port_id; // @[XConverter.scala 61:33]
  wire  fifo_h2c_cmd_io_out_bits_no_dma; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_in_clk; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_clk; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_rstn; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_in_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_in_valid; // @[XConverter.scala 61:33]
  wire [63:0] fifo_c2h_cmd_io_in_bits_addr; // @[XConverter.scala 61:33]
  wire [10:0] fifo_c2h_cmd_io_in_bits_qid; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_in_bits_error; // @[XConverter.scala 61:33]
  wire [7:0] fifo_c2h_cmd_io_in_bits_func; // @[XConverter.scala 61:33]
  wire [2:0] fifo_c2h_cmd_io_in_bits_port_id; // @[XConverter.scala 61:33]
  wire [6:0] fifo_c2h_cmd_io_in_bits_pfch_tag; // @[XConverter.scala 61:33]
  wire [31:0] fifo_c2h_cmd_io_in_bits_len; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_ready; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_valid; // @[XConverter.scala 61:33]
  wire [63:0] fifo_c2h_cmd_io_out_bits_addr; // @[XConverter.scala 61:33]
  wire [10:0] fifo_c2h_cmd_io_out_bits_qid; // @[XConverter.scala 61:33]
  wire  fifo_c2h_cmd_io_out_bits_error; // @[XConverter.scala 61:33]
  wire [7:0] fifo_c2h_cmd_io_out_bits_func; // @[XConverter.scala 61:33]
  wire [2:0] fifo_c2h_cmd_io_out_bits_port_id; // @[XConverter.scala 61:33]
  wire [6:0] fifo_c2h_cmd_io_out_bits_pfch_tag; // @[XConverter.scala 61:33]
  wire  check_c2h_clock; // @[QDMA.scala 84:95]
  wire  check_c2h_reset; // @[QDMA.scala 84:95]
  wire  check_c2h_io_in_ready; // @[QDMA.scala 84:95]
  wire  check_c2h_io_in_valid; // @[QDMA.scala 84:95]
  wire [63:0] check_c2h_io_in_bits_addr; // @[QDMA.scala 84:95]
  wire [6:0] check_c2h_io_in_bits_pfch_tag; // @[QDMA.scala 84:95]
  wire [31:0] check_c2h_io_in_bits_len; // @[QDMA.scala 84:95]
  wire  check_c2h_io_out_ready; // @[QDMA.scala 84:95]
  wire  check_c2h_io_out_valid; // @[QDMA.scala 84:95]
  wire [63:0] check_c2h_io_out_bits_addr; // @[QDMA.scala 84:95]
  wire [6:0] check_c2h_io_out_bits_pfch_tag; // @[QDMA.scala 84:95]
  wire [31:0] check_c2h_io_out_bits_len; // @[QDMA.scala 84:95]
  wire  check_h2c_clock; // @[QDMA.scala 86:95]
  wire  check_h2c_reset; // @[QDMA.scala 86:95]
  wire  check_h2c_io_in_ready; // @[QDMA.scala 86:95]
  wire  check_h2c_io_in_valid; // @[QDMA.scala 86:95]
  wire [63:0] check_h2c_io_in_bits_addr; // @[QDMA.scala 86:95]
  wire [31:0] check_h2c_io_in_bits_len; // @[QDMA.scala 86:95]
  wire  check_h2c_io_out_ready; // @[QDMA.scala 86:95]
  wire  check_h2c_io_out_valid; // @[QDMA.scala 86:95]
  wire [63:0] check_h2c_io_out_bits_addr; // @[QDMA.scala 86:95]
  wire [31:0] check_h2c_io_out_bits_len; // @[QDMA.scala 86:95]
  wire  check_h2c_io_out_bits_eop; // @[QDMA.scala 86:95]
  wire  check_h2c_io_out_bits_sop; // @[QDMA.scala 86:95]
  wire  tlb_clock; // @[QDMA.scala 89:87]
  wire  tlb_reset; // @[QDMA.scala 89:87]
  wire  tlb_io_wr_tlb_ready; // @[QDMA.scala 89:87]
  wire  tlb_io_wr_tlb_valid; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_wr_tlb_bits_vaddr_high; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_wr_tlb_bits_vaddr_low; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_wr_tlb_bits_paddr_high; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_wr_tlb_bits_paddr_low; // @[QDMA.scala 89:87]
  wire  tlb_io_wr_tlb_bits_is_base; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_in_ready; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_in_valid; // @[QDMA.scala 89:87]
  wire [63:0] tlb_io_h2c_in_bits_addr; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_h2c_in_bits_len; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_in_bits_eop; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_in_bits_sop; // @[QDMA.scala 89:87]
  wire  tlb_io_c2h_in_ready; // @[QDMA.scala 89:87]
  wire  tlb_io_c2h_in_valid; // @[QDMA.scala 89:87]
  wire [63:0] tlb_io_c2h_in_bits_addr; // @[QDMA.scala 89:87]
  wire [6:0] tlb_io_c2h_in_bits_pfch_tag; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_c2h_in_bits_len; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_out_ready; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_out_valid; // @[QDMA.scala 89:87]
  wire [63:0] tlb_io_h2c_out_bits_addr; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_h2c_out_bits_len; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_out_bits_eop; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_out_bits_sop; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_out_bits_mrkr_req; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_out_bits_sdi; // @[QDMA.scala 89:87]
  wire [10:0] tlb_io_h2c_out_bits_qid; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_out_bits_error; // @[QDMA.scala 89:87]
  wire [7:0] tlb_io_h2c_out_bits_func; // @[QDMA.scala 89:87]
  wire [15:0] tlb_io_h2c_out_bits_cidx; // @[QDMA.scala 89:87]
  wire [2:0] tlb_io_h2c_out_bits_port_id; // @[QDMA.scala 89:87]
  wire  tlb_io_h2c_out_bits_no_dma; // @[QDMA.scala 89:87]
  wire  tlb_io_c2h_out_ready; // @[QDMA.scala 89:87]
  wire  tlb_io_c2h_out_valid; // @[QDMA.scala 89:87]
  wire [63:0] tlb_io_c2h_out_bits_addr; // @[QDMA.scala 89:87]
  wire [10:0] tlb_io_c2h_out_bits_qid; // @[QDMA.scala 89:87]
  wire  tlb_io_c2h_out_bits_error; // @[QDMA.scala 89:87]
  wire [7:0] tlb_io_c2h_out_bits_func; // @[QDMA.scala 89:87]
  wire [2:0] tlb_io_c2h_out_bits_port_id; // @[QDMA.scala 89:87]
  wire [6:0] tlb_io_c2h_out_bits_pfch_tag; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_c2h_out_bits_len; // @[QDMA.scala 89:87]
  wire [31:0] tlb_io_tlb_miss_count; // @[QDMA.scala 89:87]
  wire  fifo_wr_tlb_io_in_clk; // @[XConverter.scala 61:33]
  wire  fifo_wr_tlb_io_out_clk; // @[XConverter.scala 61:33]
  wire  fifo_wr_tlb_io_rstn; // @[XConverter.scala 61:33]
  wire  fifo_wr_tlb_io_in_valid; // @[XConverter.scala 61:33]
  wire [31:0] fifo_wr_tlb_io_in_bits_vaddr_high; // @[XConverter.scala 61:33]
  wire [31:0] fifo_wr_tlb_io_in_bits_vaddr_low; // @[XConverter.scala 61:33]
  wire [31:0] fifo_wr_tlb_io_in_bits_paddr_high; // @[XConverter.scala 61:33]
  wire [31:0] fifo_wr_tlb_io_in_bits_paddr_low; // @[XConverter.scala 61:33]
  wire  fifo_wr_tlb_io_in_bits_is_base; // @[XConverter.scala 61:33]
  wire  fifo_wr_tlb_io_out_valid; // @[XConverter.scala 61:33]
  wire [31:0] fifo_wr_tlb_io_out_bits_vaddr_high; // @[XConverter.scala 61:33]
  wire [31:0] fifo_wr_tlb_io_out_bits_vaddr_low; // @[XConverter.scala 61:33]
  wire [31:0] fifo_wr_tlb_io_out_bits_paddr_high; // @[XConverter.scala 61:33]
  wire [31:0] fifo_wr_tlb_io_out_bits_paddr_low; // @[XConverter.scala 61:33]
  wire  fifo_wr_tlb_io_out_bits_is_base; // @[XConverter.scala 61:33]
  wire  axil2reg_clock; // @[QDMA.scala 108:76]
  wire  axil2reg_reset; // @[QDMA.scala 108:76]
  wire  axil2reg_io_axi_aw_ready; // @[QDMA.scala 108:76]
  wire  axil2reg_io_axi_aw_valid; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_axi_aw_bits_addr; // @[QDMA.scala 108:76]
  wire  axil2reg_io_axi_ar_ready; // @[QDMA.scala 108:76]
  wire  axil2reg_io_axi_ar_valid; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_axi_ar_bits_addr; // @[QDMA.scala 108:76]
  wire  axil2reg_io_axi_w_ready; // @[QDMA.scala 108:76]
  wire  axil2reg_io_axi_w_valid; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_axi_w_bits_data; // @[QDMA.scala 108:76]
  wire  axil2reg_io_axi_r_ready; // @[QDMA.scala 108:76]
  wire  axil2reg_io_axi_r_valid; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_axi_r_bits_data; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_8; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_9; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_10; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_11; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_12; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_13; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_20; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_50; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_51; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_52; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_53; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_54; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_55; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_56; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_57; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_58; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_59; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_70; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_71; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_72; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_73; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_74; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_75; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_76; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_77; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_78; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_79; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_80; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_91; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_92; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_93; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_control_94; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_40; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_51; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_52; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_61; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_71; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_72; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_75; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_76; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_77; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_78; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_79; // @[QDMA.scala 108:76]
  wire [31:0] axil2reg_io_reg_status_81; // @[QDMA.scala 108:76]
  wire  boundary_split_clock; // @[QDMA.scala 126:103]
  wire  boundary_split_reset; // @[QDMA.scala 126:103]
  wire  boundary_split_io_data_in_ready; // @[QDMA.scala 126:103]
  wire  boundary_split_io_data_in_valid; // @[QDMA.scala 126:103]
  wire [511:0] boundary_split_io_data_in_bits_data; // @[QDMA.scala 126:103]
  wire  boundary_split_io_cmd_in_ready; // @[QDMA.scala 126:103]
  wire  boundary_split_io_cmd_in_valid; // @[QDMA.scala 126:103]
  wire [63:0] boundary_split_io_cmd_in_bits_addr; // @[QDMA.scala 126:103]
  wire [10:0] boundary_split_io_cmd_in_bits_qid; // @[QDMA.scala 126:103]
  wire  boundary_split_io_cmd_in_bits_error; // @[QDMA.scala 126:103]
  wire [7:0] boundary_split_io_cmd_in_bits_func; // @[QDMA.scala 126:103]
  wire [2:0] boundary_split_io_cmd_in_bits_port_id; // @[QDMA.scala 126:103]
  wire [6:0] boundary_split_io_cmd_in_bits_pfch_tag; // @[QDMA.scala 126:103]
  wire [31:0] boundary_split_io_cmd_in_bits_len; // @[QDMA.scala 126:103]
  wire  boundary_split_io_data_out_ready; // @[QDMA.scala 126:103]
  wire  boundary_split_io_data_out_valid; // @[QDMA.scala 126:103]
  wire [511:0] boundary_split_io_data_out_bits_data; // @[QDMA.scala 126:103]
  wire [31:0] boundary_split_io_data_out_bits_tcrc; // @[QDMA.scala 126:103]
  wire  boundary_split_io_data_out_bits_ctrl_marker; // @[QDMA.scala 126:103]
  wire [6:0] boundary_split_io_data_out_bits_ctrl_ecc; // @[QDMA.scala 126:103]
  wire [31:0] boundary_split_io_data_out_bits_ctrl_len; // @[QDMA.scala 126:103]
  wire [2:0] boundary_split_io_data_out_bits_ctrl_port_id; // @[QDMA.scala 126:103]
  wire [10:0] boundary_split_io_data_out_bits_ctrl_qid; // @[QDMA.scala 126:103]
  wire  boundary_split_io_data_out_bits_ctrl_has_cmpt; // @[QDMA.scala 126:103]
  wire  boundary_split_io_data_out_bits_last; // @[QDMA.scala 126:103]
  wire [5:0] boundary_split_io_data_out_bits_mty; // @[QDMA.scala 126:103]
  wire  boundary_split_io_cmd_out_ready; // @[QDMA.scala 126:103]
  wire  boundary_split_io_cmd_out_valid; // @[QDMA.scala 126:103]
  wire [63:0] boundary_split_io_cmd_out_bits_addr; // @[QDMA.scala 126:103]
  wire [10:0] boundary_split_io_cmd_out_bits_qid; // @[QDMA.scala 126:103]
  wire  boundary_split_io_cmd_out_bits_error; // @[QDMA.scala 126:103]
  wire [7:0] boundary_split_io_cmd_out_bits_func; // @[QDMA.scala 126:103]
  wire [2:0] boundary_split_io_cmd_out_bits_port_id; // @[QDMA.scala 126:103]
  wire [6:0] boundary_split_io_cmd_out_bits_pfch_tag; // @[QDMA.scala 126:103]
  wire [31:0] boundary_split_io_cmd_out_bits_len; // @[QDMA.scala 126:103]
  wire  qdma_inst_sys_rst_n; // @[QDMA.scala 133:31]
  wire  qdma_inst_sys_clk; // @[QDMA.scala 133:31]
  wire  qdma_inst_sys_clk_gt; // @[QDMA.scala 133:31]
  wire [15:0] qdma_inst_pci_exp_txn; // @[QDMA.scala 133:31]
  wire [15:0] qdma_inst_pci_exp_txp; // @[QDMA.scala 133:31]
  wire [15:0] qdma_inst_pci_exp_rxn; // @[QDMA.scala 133:31]
  wire [15:0] qdma_inst_pci_exp_rxp; // @[QDMA.scala 133:31]
  wire [3:0] qdma_inst_m_axib_awid; // @[QDMA.scala 133:31]
  wire [63:0] qdma_inst_m_axib_awaddr; // @[QDMA.scala 133:31]
  wire [7:0] qdma_inst_m_axib_awlen; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_m_axib_awsize; // @[QDMA.scala 133:31]
  wire [1:0] qdma_inst_m_axib_awburst; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_m_axib_awprot; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_awlock; // @[QDMA.scala 133:31]
  wire [3:0] qdma_inst_m_axib_awcache; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_awvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_awready; // @[QDMA.scala 133:31]
  wire [511:0] qdma_inst_m_axib_wdata; // @[QDMA.scala 133:31]
  wire [63:0] qdma_inst_m_axib_wstrb; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_wlast; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_wvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_wready; // @[QDMA.scala 133:31]
  wire [3:0] qdma_inst_m_axib_bid; // @[QDMA.scala 133:31]
  wire [1:0] qdma_inst_m_axib_bresp; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_bvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_bready; // @[QDMA.scala 133:31]
  wire [3:0] qdma_inst_m_axib_arid; // @[QDMA.scala 133:31]
  wire [63:0] qdma_inst_m_axib_araddr; // @[QDMA.scala 133:31]
  wire [7:0] qdma_inst_m_axib_arlen; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_m_axib_arsize; // @[QDMA.scala 133:31]
  wire [1:0] qdma_inst_m_axib_arburst; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_m_axib_arprot; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_arlock; // @[QDMA.scala 133:31]
  wire [3:0] qdma_inst_m_axib_arcache; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_arvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_arready; // @[QDMA.scala 133:31]
  wire [3:0] qdma_inst_m_axib_rid; // @[QDMA.scala 133:31]
  wire [511:0] qdma_inst_m_axib_rdata; // @[QDMA.scala 133:31]
  wire [1:0] qdma_inst_m_axib_rresp; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_rlast; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_rvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axib_rready; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_m_axil_awaddr; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_awvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_awready; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_m_axil_wdata; // @[QDMA.scala 133:31]
  wire [3:0] qdma_inst_m_axil_wstrb; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_wvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_wready; // @[QDMA.scala 133:31]
  wire [1:0] qdma_inst_m_axil_bresp; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_bvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_bready; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_m_axil_araddr; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_arvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_arready; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_m_axil_rdata; // @[QDMA.scala 133:31]
  wire [1:0] qdma_inst_m_axil_rresp; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_rvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axil_rready; // @[QDMA.scala 133:31]
  wire  qdma_inst_axi_aclk; // @[QDMA.scala 133:31]
  wire  qdma_inst_axi_aresetn; // @[QDMA.scala 133:31]
  wire  qdma_inst_soft_reset_n; // @[QDMA.scala 133:31]
  wire [63:0] qdma_inst_h2c_byp_in_st_addr; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_h2c_byp_in_st_len; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_in_st_eop; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_in_st_sop; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_in_st_mrkr_req; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_in_st_sdi; // @[QDMA.scala 133:31]
  wire [10:0] qdma_inst_h2c_byp_in_st_qid; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_in_st_error; // @[QDMA.scala 133:31]
  wire [7:0] qdma_inst_h2c_byp_in_st_func; // @[QDMA.scala 133:31]
  wire [15:0] qdma_inst_h2c_byp_in_st_cidx; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_h2c_byp_in_st_port_id; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_in_st_no_dma; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_in_st_vld; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_in_st_rdy; // @[QDMA.scala 133:31]
  wire [63:0] qdma_inst_c2h_byp_in_st_csh_addr; // @[QDMA.scala 133:31]
  wire [10:0] qdma_inst_c2h_byp_in_st_csh_qid; // @[QDMA.scala 133:31]
  wire  qdma_inst_c2h_byp_in_st_csh_error; // @[QDMA.scala 133:31]
  wire [7:0] qdma_inst_c2h_byp_in_st_csh_func; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_c2h_byp_in_st_csh_port_id; // @[QDMA.scala 133:31]
  wire [6:0] qdma_inst_c2h_byp_in_st_csh_pfch_tag; // @[QDMA.scala 133:31]
  wire  qdma_inst_c2h_byp_in_st_csh_vld; // @[QDMA.scala 133:31]
  wire  qdma_inst_c2h_byp_in_st_csh_rdy; // @[QDMA.scala 133:31]
  wire [511:0] qdma_inst_s_axis_c2h_tdata; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_s_axis_c2h_tcrc; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_ctrl_marker; // @[QDMA.scala 133:31]
  wire [6:0] qdma_inst_s_axis_c2h_ctrl_ecc; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_s_axis_c2h_ctrl_len; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_s_axis_c2h_ctrl_port_id; // @[QDMA.scala 133:31]
  wire [10:0] qdma_inst_s_axis_c2h_ctrl_qid; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_ctrl_has_cmpt; // @[QDMA.scala 133:31]
  wire [5:0] qdma_inst_s_axis_c2h_mty; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_tlast; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_tvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_tready; // @[QDMA.scala 133:31]
  wire [511:0] qdma_inst_m_axis_h2c_tdata; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_m_axis_h2c_tcrc; // @[QDMA.scala 133:31]
  wire [10:0] qdma_inst_m_axis_h2c_tuser_qid; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_m_axis_h2c_tuser_port_id; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axis_h2c_tuser_err; // @[QDMA.scala 133:31]
  wire [31:0] qdma_inst_m_axis_h2c_tuser_mdata; // @[QDMA.scala 133:31]
  wire [5:0] qdma_inst_m_axis_h2c_tuser_mty; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axis_h2c_tuser_zero_byte; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axis_h2c_tlast; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axis_h2c_tvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_m_axis_h2c_tready; // @[QDMA.scala 133:31]
  wire  qdma_inst_axis_c2h_status_drop; // @[QDMA.scala 133:31]
  wire  qdma_inst_axis_c2h_status_last; // @[QDMA.scala 133:31]
  wire  qdma_inst_axis_c2h_status_cmp; // @[QDMA.scala 133:31]
  wire  qdma_inst_axis_c2h_status_valid; // @[QDMA.scala 133:31]
  wire  qdma_inst_axis_c2h_status_error; // @[QDMA.scala 133:31]
  wire [10:0] qdma_inst_axis_c2h_status_qid; // @[QDMA.scala 133:31]
  wire [511:0] qdma_inst_s_axis_c2h_cmpt_tdata; // @[QDMA.scala 133:31]
  wire [1:0] qdma_inst_s_axis_c2h_cmpt_size; // @[QDMA.scala 133:31]
  wire [15:0] qdma_inst_s_axis_c2h_cmpt_dpar; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_cmpt_tvalid; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_cmpt_tready; // @[QDMA.scala 133:31]
  wire [10:0] qdma_inst_s_axis_c2h_cmpt_ctrl_qid; // @[QDMA.scala 133:31]
  wire [1:0] qdma_inst_s_axis_c2h_cmpt_ctrl_cmpt_type; // @[QDMA.scala 133:31]
  wire [15:0] qdma_inst_s_axis_c2h_cmpt_ctrl_wait_pld_pkt_id; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_cmpt_ctrl_no_wrb_marker; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_s_axis_c2h_cmpt_ctrl_port_id; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_cmpt_ctrl_marker; // @[QDMA.scala 133:31]
  wire  qdma_inst_s_axis_c2h_cmpt_ctrl_user_trig; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_s_axis_c2h_cmpt_ctrl_col_idx; // @[QDMA.scala 133:31]
  wire [2:0] qdma_inst_s_axis_c2h_cmpt_ctrl_err_idx; // @[QDMA.scala 133:31]
  wire  qdma_inst_h2c_byp_out_rdy; // @[QDMA.scala 133:31]
  wire  qdma_inst_c2h_byp_out_rdy; // @[QDMA.scala 133:31]
  wire  qdma_inst_tm_dsc_sts_rdy; // @[QDMA.scala 133:31]
  wire  qdma_inst_dsc_crdt_in_vld; // @[QDMA.scala 133:31]
  wire  qdma_inst_dsc_crdt_in_rdy; // @[QDMA.scala 133:31]
  wire  qdma_inst_dsc_crdt_in_dir; // @[QDMA.scala 133:31]
  wire  qdma_inst_dsc_crdt_in_fence; // @[QDMA.scala 133:31]
  wire [10:0] qdma_inst_dsc_crdt_in_qid; // @[QDMA.scala 133:31]
  wire [15:0] qdma_inst_dsc_crdt_in_crdt; // @[QDMA.scala 133:31]
  wire  qdma_inst_qsts_out_rdy; // @[QDMA.scala 133:31]
  wire  qdma_inst_usr_irq_in_vld; // @[QDMA.scala 133:31]
  wire [10:0] qdma_inst_usr_irq_in_vec; // @[QDMA.scala 133:31]
  wire [7:0] qdma_inst_usr_irq_in_fnc; // @[QDMA.scala 133:31]
  wire  qdma_inst_usr_irq_out_ack; // @[QDMA.scala 133:31]
  wire  qdma_inst_usr_irq_out_fail; // @[QDMA.scala 133:31]
  reg  fifo_wr_tlb_io_in_valid_REG; // @[QDMA.scala 102:107]
  reg  fifo_wr_tlb_io_in_valid_REG_1; // @[QDMA.scala 102:98]
  IBUF perst_n_pad ( // @[Buf.scala 17:34]
    .O(perst_n_pad_O),
    .I(perst_n_pad_I)
  );
  IBUFDS_GTE4 #(.REFCLK_EN_TX_PATH(0), .REFCLK_HROW_CK_SEL(0), .REFCLK_ICNTL_RX(0)) ibufds_gte4_inst ( // @[QDMA.scala 70:38]
    .O(ibufds_gte4_inst_O),
    .ODIV2(ibufds_gte4_inst_ODIV2),
    .CEB(ibufds_gte4_inst_CEB),
    .I(ibufds_gte4_inst_I),
    .IB(ibufds_gte4_inst_IB)
  );
  XConverter fifo_h2c_data ( // @[XConverter.scala 61:33]
    .io_in_clk(fifo_h2c_data_io_in_clk),
    .io_out_clk(fifo_h2c_data_io_out_clk),
    .io_rstn(fifo_h2c_data_io_rstn),
    .io_in_ready(fifo_h2c_data_io_in_ready),
    .io_in_valid(fifo_h2c_data_io_in_valid),
    .io_in_bits_data(fifo_h2c_data_io_in_bits_data),
    .io_in_bits_tcrc(fifo_h2c_data_io_in_bits_tcrc),
    .io_in_bits_tuser_qid(fifo_h2c_data_io_in_bits_tuser_qid),
    .io_in_bits_tuser_port_id(fifo_h2c_data_io_in_bits_tuser_port_id),
    .io_in_bits_tuser_err(fifo_h2c_data_io_in_bits_tuser_err),
    .io_in_bits_tuser_mdata(fifo_h2c_data_io_in_bits_tuser_mdata),
    .io_in_bits_tuser_mty(fifo_h2c_data_io_in_bits_tuser_mty),
    .io_in_bits_tuser_zero_byte(fifo_h2c_data_io_in_bits_tuser_zero_byte),
    .io_in_bits_last(fifo_h2c_data_io_in_bits_last),
    .io_out_ready(fifo_h2c_data_io_out_ready),
    .io_out_valid(fifo_h2c_data_io_out_valid),
    .io_out_bits_data(fifo_h2c_data_io_out_bits_data)
  );
  XConverter_1 fifo_c2h_data ( // @[XConverter.scala 61:33]
    .io_in_clk(fifo_c2h_data_io_in_clk),
    .io_out_clk(fifo_c2h_data_io_out_clk),
    .io_rstn(fifo_c2h_data_io_rstn),
    .io_in_ready(fifo_c2h_data_io_in_ready),
    .io_in_valid(fifo_c2h_data_io_in_valid),
    .io_in_bits_data(fifo_c2h_data_io_in_bits_data),
    .io_in_bits_tcrc(fifo_c2h_data_io_in_bits_tcrc),
    .io_in_bits_ctrl_marker(fifo_c2h_data_io_in_bits_ctrl_marker),
    .io_in_bits_ctrl_ecc(fifo_c2h_data_io_in_bits_ctrl_ecc),
    .io_in_bits_ctrl_len(fifo_c2h_data_io_in_bits_ctrl_len),
    .io_in_bits_ctrl_port_id(fifo_c2h_data_io_in_bits_ctrl_port_id),
    .io_in_bits_ctrl_qid(fifo_c2h_data_io_in_bits_ctrl_qid),
    .io_in_bits_ctrl_has_cmpt(fifo_c2h_data_io_in_bits_ctrl_has_cmpt),
    .io_in_bits_last(fifo_c2h_data_io_in_bits_last),
    .io_in_bits_mty(fifo_c2h_data_io_in_bits_mty),
    .io_out_ready(fifo_c2h_data_io_out_ready),
    .io_out_valid(fifo_c2h_data_io_out_valid),
    .io_out_bits_data(fifo_c2h_data_io_out_bits_data),
    .io_out_bits_tcrc(fifo_c2h_data_io_out_bits_tcrc),
    .io_out_bits_ctrl_marker(fifo_c2h_data_io_out_bits_ctrl_marker),
    .io_out_bits_ctrl_ecc(fifo_c2h_data_io_out_bits_ctrl_ecc),
    .io_out_bits_ctrl_len(fifo_c2h_data_io_out_bits_ctrl_len),
    .io_out_bits_ctrl_port_id(fifo_c2h_data_io_out_bits_ctrl_port_id),
    .io_out_bits_ctrl_qid(fifo_c2h_data_io_out_bits_ctrl_qid),
    .io_out_bits_ctrl_has_cmpt(fifo_c2h_data_io_out_bits_ctrl_has_cmpt),
    .io_out_bits_last(fifo_c2h_data_io_out_bits_last),
    .io_out_bits_mty(fifo_c2h_data_io_out_bits_mty)
  );
  XConverter_2 fifo_h2c_cmd ( // @[XConverter.scala 61:33]
    .io_in_clk(fifo_h2c_cmd_io_in_clk),
    .io_out_clk(fifo_h2c_cmd_io_out_clk),
    .io_rstn(fifo_h2c_cmd_io_rstn),
    .io_in_ready(fifo_h2c_cmd_io_in_ready),
    .io_in_valid(fifo_h2c_cmd_io_in_valid),
    .io_in_bits_addr(fifo_h2c_cmd_io_in_bits_addr),
    .io_in_bits_len(fifo_h2c_cmd_io_in_bits_len),
    .io_in_bits_eop(fifo_h2c_cmd_io_in_bits_eop),
    .io_in_bits_sop(fifo_h2c_cmd_io_in_bits_sop),
    .io_in_bits_mrkr_req(fifo_h2c_cmd_io_in_bits_mrkr_req),
    .io_in_bits_sdi(fifo_h2c_cmd_io_in_bits_sdi),
    .io_in_bits_qid(fifo_h2c_cmd_io_in_bits_qid),
    .io_in_bits_error(fifo_h2c_cmd_io_in_bits_error),
    .io_in_bits_func(fifo_h2c_cmd_io_in_bits_func),
    .io_in_bits_cidx(fifo_h2c_cmd_io_in_bits_cidx),
    .io_in_bits_port_id(fifo_h2c_cmd_io_in_bits_port_id),
    .io_in_bits_no_dma(fifo_h2c_cmd_io_in_bits_no_dma),
    .io_out_ready(fifo_h2c_cmd_io_out_ready),
    .io_out_valid(fifo_h2c_cmd_io_out_valid),
    .io_out_bits_addr(fifo_h2c_cmd_io_out_bits_addr),
    .io_out_bits_len(fifo_h2c_cmd_io_out_bits_len),
    .io_out_bits_eop(fifo_h2c_cmd_io_out_bits_eop),
    .io_out_bits_sop(fifo_h2c_cmd_io_out_bits_sop),
    .io_out_bits_mrkr_req(fifo_h2c_cmd_io_out_bits_mrkr_req),
    .io_out_bits_sdi(fifo_h2c_cmd_io_out_bits_sdi),
    .io_out_bits_qid(fifo_h2c_cmd_io_out_bits_qid),
    .io_out_bits_error(fifo_h2c_cmd_io_out_bits_error),
    .io_out_bits_func(fifo_h2c_cmd_io_out_bits_func),
    .io_out_bits_cidx(fifo_h2c_cmd_io_out_bits_cidx),
    .io_out_bits_port_id(fifo_h2c_cmd_io_out_bits_port_id),
    .io_out_bits_no_dma(fifo_h2c_cmd_io_out_bits_no_dma)
  );
  XConverter_3 fifo_c2h_cmd ( // @[XConverter.scala 61:33]
    .io_in_clk(fifo_c2h_cmd_io_in_clk),
    .io_out_clk(fifo_c2h_cmd_io_out_clk),
    .io_rstn(fifo_c2h_cmd_io_rstn),
    .io_in_ready(fifo_c2h_cmd_io_in_ready),
    .io_in_valid(fifo_c2h_cmd_io_in_valid),
    .io_in_bits_addr(fifo_c2h_cmd_io_in_bits_addr),
    .io_in_bits_qid(fifo_c2h_cmd_io_in_bits_qid),
    .io_in_bits_error(fifo_c2h_cmd_io_in_bits_error),
    .io_in_bits_func(fifo_c2h_cmd_io_in_bits_func),
    .io_in_bits_port_id(fifo_c2h_cmd_io_in_bits_port_id),
    .io_in_bits_pfch_tag(fifo_c2h_cmd_io_in_bits_pfch_tag),
    .io_in_bits_len(fifo_c2h_cmd_io_in_bits_len),
    .io_out_ready(fifo_c2h_cmd_io_out_ready),
    .io_out_valid(fifo_c2h_cmd_io_out_valid),
    .io_out_bits_addr(fifo_c2h_cmd_io_out_bits_addr),
    .io_out_bits_qid(fifo_c2h_cmd_io_out_bits_qid),
    .io_out_bits_error(fifo_c2h_cmd_io_out_bits_error),
    .io_out_bits_func(fifo_c2h_cmd_io_out_bits_func),
    .io_out_bits_port_id(fifo_c2h_cmd_io_out_bits_port_id),
    .io_out_bits_pfch_tag(fifo_c2h_cmd_io_out_bits_pfch_tag)
  );
  CMDBoundaryCheck check_c2h ( // @[QDMA.scala 84:95]
    .clock(check_c2h_clock),
    .reset(check_c2h_reset),
    .io_in_ready(check_c2h_io_in_ready),
    .io_in_valid(check_c2h_io_in_valid),
    .io_in_bits_addr(check_c2h_io_in_bits_addr),
    .io_in_bits_pfch_tag(check_c2h_io_in_bits_pfch_tag),
    .io_in_bits_len(check_c2h_io_in_bits_len),
    .io_out_ready(check_c2h_io_out_ready),
    .io_out_valid(check_c2h_io_out_valid),
    .io_out_bits_addr(check_c2h_io_out_bits_addr),
    .io_out_bits_pfch_tag(check_c2h_io_out_bits_pfch_tag),
    .io_out_bits_len(check_c2h_io_out_bits_len)
  );
  CMDBoundaryCheck_1 check_h2c ( // @[QDMA.scala 86:95]
    .clock(check_h2c_clock),
    .reset(check_h2c_reset),
    .io_in_ready(check_h2c_io_in_ready),
    .io_in_valid(check_h2c_io_in_valid),
    .io_in_bits_addr(check_h2c_io_in_bits_addr),
    .io_in_bits_len(check_h2c_io_in_bits_len),
    .io_out_ready(check_h2c_io_out_ready),
    .io_out_valid(check_h2c_io_out_valid),
    .io_out_bits_addr(check_h2c_io_out_bits_addr),
    .io_out_bits_len(check_h2c_io_out_bits_len),
    .io_out_bits_eop(check_h2c_io_out_bits_eop),
    .io_out_bits_sop(check_h2c_io_out_bits_sop)
  );
  TLB tlb ( // @[QDMA.scala 89:87]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_wr_tlb_ready(tlb_io_wr_tlb_ready),
    .io_wr_tlb_valid(tlb_io_wr_tlb_valid),
    .io_wr_tlb_bits_vaddr_high(tlb_io_wr_tlb_bits_vaddr_high),
    .io_wr_tlb_bits_vaddr_low(tlb_io_wr_tlb_bits_vaddr_low),
    .io_wr_tlb_bits_paddr_high(tlb_io_wr_tlb_bits_paddr_high),
    .io_wr_tlb_bits_paddr_low(tlb_io_wr_tlb_bits_paddr_low),
    .io_wr_tlb_bits_is_base(tlb_io_wr_tlb_bits_is_base),
    .io_h2c_in_ready(tlb_io_h2c_in_ready),
    .io_h2c_in_valid(tlb_io_h2c_in_valid),
    .io_h2c_in_bits_addr(tlb_io_h2c_in_bits_addr),
    .io_h2c_in_bits_len(tlb_io_h2c_in_bits_len),
    .io_h2c_in_bits_eop(tlb_io_h2c_in_bits_eop),
    .io_h2c_in_bits_sop(tlb_io_h2c_in_bits_sop),
    .io_c2h_in_ready(tlb_io_c2h_in_ready),
    .io_c2h_in_valid(tlb_io_c2h_in_valid),
    .io_c2h_in_bits_addr(tlb_io_c2h_in_bits_addr),
    .io_c2h_in_bits_pfch_tag(tlb_io_c2h_in_bits_pfch_tag),
    .io_c2h_in_bits_len(tlb_io_c2h_in_bits_len),
    .io_h2c_out_ready(tlb_io_h2c_out_ready),
    .io_h2c_out_valid(tlb_io_h2c_out_valid),
    .io_h2c_out_bits_addr(tlb_io_h2c_out_bits_addr),
    .io_h2c_out_bits_len(tlb_io_h2c_out_bits_len),
    .io_h2c_out_bits_eop(tlb_io_h2c_out_bits_eop),
    .io_h2c_out_bits_sop(tlb_io_h2c_out_bits_sop),
    .io_h2c_out_bits_mrkr_req(tlb_io_h2c_out_bits_mrkr_req),
    .io_h2c_out_bits_sdi(tlb_io_h2c_out_bits_sdi),
    .io_h2c_out_bits_qid(tlb_io_h2c_out_bits_qid),
    .io_h2c_out_bits_error(tlb_io_h2c_out_bits_error),
    .io_h2c_out_bits_func(tlb_io_h2c_out_bits_func),
    .io_h2c_out_bits_cidx(tlb_io_h2c_out_bits_cidx),
    .io_h2c_out_bits_port_id(tlb_io_h2c_out_bits_port_id),
    .io_h2c_out_bits_no_dma(tlb_io_h2c_out_bits_no_dma),
    .io_c2h_out_ready(tlb_io_c2h_out_ready),
    .io_c2h_out_valid(tlb_io_c2h_out_valid),
    .io_c2h_out_bits_addr(tlb_io_c2h_out_bits_addr),
    .io_c2h_out_bits_qid(tlb_io_c2h_out_bits_qid),
    .io_c2h_out_bits_error(tlb_io_c2h_out_bits_error),
    .io_c2h_out_bits_func(tlb_io_c2h_out_bits_func),
    .io_c2h_out_bits_port_id(tlb_io_c2h_out_bits_port_id),
    .io_c2h_out_bits_pfch_tag(tlb_io_c2h_out_bits_pfch_tag),
    .io_c2h_out_bits_len(tlb_io_c2h_out_bits_len),
    .io_tlb_miss_count(tlb_io_tlb_miss_count)
  );
  XConverter_4 fifo_wr_tlb ( // @[XConverter.scala 61:33]
    .io_in_clk(fifo_wr_tlb_io_in_clk),
    .io_out_clk(fifo_wr_tlb_io_out_clk),
    .io_rstn(fifo_wr_tlb_io_rstn),
    .io_in_valid(fifo_wr_tlb_io_in_valid),
    .io_in_bits_vaddr_high(fifo_wr_tlb_io_in_bits_vaddr_high),
    .io_in_bits_vaddr_low(fifo_wr_tlb_io_in_bits_vaddr_low),
    .io_in_bits_paddr_high(fifo_wr_tlb_io_in_bits_paddr_high),
    .io_in_bits_paddr_low(fifo_wr_tlb_io_in_bits_paddr_low),
    .io_in_bits_is_base(fifo_wr_tlb_io_in_bits_is_base),
    .io_out_valid(fifo_wr_tlb_io_out_valid),
    .io_out_bits_vaddr_high(fifo_wr_tlb_io_out_bits_vaddr_high),
    .io_out_bits_vaddr_low(fifo_wr_tlb_io_out_bits_vaddr_low),
    .io_out_bits_paddr_high(fifo_wr_tlb_io_out_bits_paddr_high),
    .io_out_bits_paddr_low(fifo_wr_tlb_io_out_bits_paddr_low),
    .io_out_bits_is_base(fifo_wr_tlb_io_out_bits_is_base)
  );
  PoorAXIL2Reg axil2reg ( // @[QDMA.scala 108:76]
    .clock(axil2reg_clock),
    .reset(axil2reg_reset),
    .io_axi_aw_ready(axil2reg_io_axi_aw_ready),
    .io_axi_aw_valid(axil2reg_io_axi_aw_valid),
    .io_axi_aw_bits_addr(axil2reg_io_axi_aw_bits_addr),
    .io_axi_ar_ready(axil2reg_io_axi_ar_ready),
    .io_axi_ar_valid(axil2reg_io_axi_ar_valid),
    .io_axi_ar_bits_addr(axil2reg_io_axi_ar_bits_addr),
    .io_axi_w_ready(axil2reg_io_axi_w_ready),
    .io_axi_w_valid(axil2reg_io_axi_w_valid),
    .io_axi_w_bits_data(axil2reg_io_axi_w_bits_data),
    .io_axi_r_ready(axil2reg_io_axi_r_ready),
    .io_axi_r_valid(axil2reg_io_axi_r_valid),
    .io_axi_r_bits_data(axil2reg_io_axi_r_bits_data),
    .io_reg_control_8(axil2reg_io_reg_control_8),
    .io_reg_control_9(axil2reg_io_reg_control_9),
    .io_reg_control_10(axil2reg_io_reg_control_10),
    .io_reg_control_11(axil2reg_io_reg_control_11),
    .io_reg_control_12(axil2reg_io_reg_control_12),
    .io_reg_control_13(axil2reg_io_reg_control_13),
    .io_reg_control_20(axil2reg_io_reg_control_20),
    .io_reg_control_50(axil2reg_io_reg_control_50),
    .io_reg_control_51(axil2reg_io_reg_control_51),
    .io_reg_control_52(axil2reg_io_reg_control_52),
    .io_reg_control_53(axil2reg_io_reg_control_53),
    .io_reg_control_54(axil2reg_io_reg_control_54),
    .io_reg_control_55(axil2reg_io_reg_control_55),
    .io_reg_control_56(axil2reg_io_reg_control_56),
    .io_reg_control_57(axil2reg_io_reg_control_57),
    .io_reg_control_58(axil2reg_io_reg_control_58),
    .io_reg_control_59(axil2reg_io_reg_control_59),
    .io_reg_control_70(axil2reg_io_reg_control_70),
    .io_reg_control_71(axil2reg_io_reg_control_71),
    .io_reg_control_72(axil2reg_io_reg_control_72),
    .io_reg_control_73(axil2reg_io_reg_control_73),
    .io_reg_control_74(axil2reg_io_reg_control_74),
    .io_reg_control_75(axil2reg_io_reg_control_75),
    .io_reg_control_76(axil2reg_io_reg_control_76),
    .io_reg_control_77(axil2reg_io_reg_control_77),
    .io_reg_control_78(axil2reg_io_reg_control_78),
    .io_reg_control_79(axil2reg_io_reg_control_79),
    .io_reg_control_80(axil2reg_io_reg_control_80),
    .io_reg_control_91(axil2reg_io_reg_control_91),
    .io_reg_control_92(axil2reg_io_reg_control_92),
    .io_reg_control_93(axil2reg_io_reg_control_93),
    .io_reg_control_94(axil2reg_io_reg_control_94),
    .io_reg_status_40(axil2reg_io_reg_status_40),
    .io_reg_status_51(axil2reg_io_reg_status_51),
    .io_reg_status_52(axil2reg_io_reg_status_52),
    .io_reg_status_61(axil2reg_io_reg_status_61),
    .io_reg_status_71(axil2reg_io_reg_status_71),
    .io_reg_status_72(axil2reg_io_reg_status_72),
    .io_reg_status_75(axil2reg_io_reg_status_75),
    .io_reg_status_76(axil2reg_io_reg_status_76),
    .io_reg_status_77(axil2reg_io_reg_status_77),
    .io_reg_status_78(axil2reg_io_reg_status_78),
    .io_reg_status_79(axil2reg_io_reg_status_79),
    .io_reg_status_81(axil2reg_io_reg_status_81)
  );
  DataBoundarySplit boundary_split ( // @[QDMA.scala 126:103]
    .clock(boundary_split_clock),
    .reset(boundary_split_reset),
    .io_data_in_ready(boundary_split_io_data_in_ready),
    .io_data_in_valid(boundary_split_io_data_in_valid),
    .io_data_in_bits_data(boundary_split_io_data_in_bits_data),
    .io_cmd_in_ready(boundary_split_io_cmd_in_ready),
    .io_cmd_in_valid(boundary_split_io_cmd_in_valid),
    .io_cmd_in_bits_addr(boundary_split_io_cmd_in_bits_addr),
    .io_cmd_in_bits_qid(boundary_split_io_cmd_in_bits_qid),
    .io_cmd_in_bits_error(boundary_split_io_cmd_in_bits_error),
    .io_cmd_in_bits_func(boundary_split_io_cmd_in_bits_func),
    .io_cmd_in_bits_port_id(boundary_split_io_cmd_in_bits_port_id),
    .io_cmd_in_bits_pfch_tag(boundary_split_io_cmd_in_bits_pfch_tag),
    .io_cmd_in_bits_len(boundary_split_io_cmd_in_bits_len),
    .io_data_out_ready(boundary_split_io_data_out_ready),
    .io_data_out_valid(boundary_split_io_data_out_valid),
    .io_data_out_bits_data(boundary_split_io_data_out_bits_data),
    .io_data_out_bits_tcrc(boundary_split_io_data_out_bits_tcrc),
    .io_data_out_bits_ctrl_marker(boundary_split_io_data_out_bits_ctrl_marker),
    .io_data_out_bits_ctrl_ecc(boundary_split_io_data_out_bits_ctrl_ecc),
    .io_data_out_bits_ctrl_len(boundary_split_io_data_out_bits_ctrl_len),
    .io_data_out_bits_ctrl_port_id(boundary_split_io_data_out_bits_ctrl_port_id),
    .io_data_out_bits_ctrl_qid(boundary_split_io_data_out_bits_ctrl_qid),
    .io_data_out_bits_ctrl_has_cmpt(boundary_split_io_data_out_bits_ctrl_has_cmpt),
    .io_data_out_bits_last(boundary_split_io_data_out_bits_last),
    .io_data_out_bits_mty(boundary_split_io_data_out_bits_mty),
    .io_cmd_out_ready(boundary_split_io_cmd_out_ready),
    .io_cmd_out_valid(boundary_split_io_cmd_out_valid),
    .io_cmd_out_bits_addr(boundary_split_io_cmd_out_bits_addr),
    .io_cmd_out_bits_qid(boundary_split_io_cmd_out_bits_qid),
    .io_cmd_out_bits_error(boundary_split_io_cmd_out_bits_error),
    .io_cmd_out_bits_func(boundary_split_io_cmd_out_bits_func),
    .io_cmd_out_bits_port_id(boundary_split_io_cmd_out_bits_port_id),
    .io_cmd_out_bits_pfch_tag(boundary_split_io_cmd_out_bits_pfch_tag),
    .io_cmd_out_bits_len(boundary_split_io_cmd_out_bits_len)
  );
  QDMABlackBox qdma_inst ( // @[QDMA.scala 133:31]
    .sys_rst_n(qdma_inst_sys_rst_n),
    .sys_clk(qdma_inst_sys_clk),
    .sys_clk_gt(qdma_inst_sys_clk_gt),
    .pci_exp_txn(qdma_inst_pci_exp_txn),
    .pci_exp_txp(qdma_inst_pci_exp_txp),
    .pci_exp_rxn(qdma_inst_pci_exp_rxn),
    .pci_exp_rxp(qdma_inst_pci_exp_rxp),
    .m_axib_awid(qdma_inst_m_axib_awid),
    .m_axib_awaddr(qdma_inst_m_axib_awaddr),
    .m_axib_awlen(qdma_inst_m_axib_awlen),
    .m_axib_awsize(qdma_inst_m_axib_awsize),
    .m_axib_awburst(qdma_inst_m_axib_awburst),
    .m_axib_awprot(qdma_inst_m_axib_awprot),
    .m_axib_awlock(qdma_inst_m_axib_awlock),
    .m_axib_awcache(qdma_inst_m_axib_awcache),
    .m_axib_awvalid(qdma_inst_m_axib_awvalid),
    .m_axib_awready(qdma_inst_m_axib_awready),
    .m_axib_wdata(qdma_inst_m_axib_wdata),
    .m_axib_wstrb(qdma_inst_m_axib_wstrb),
    .m_axib_wlast(qdma_inst_m_axib_wlast),
    .m_axib_wvalid(qdma_inst_m_axib_wvalid),
    .m_axib_wready(qdma_inst_m_axib_wready),
    .m_axib_bid(qdma_inst_m_axib_bid),
    .m_axib_bresp(qdma_inst_m_axib_bresp),
    .m_axib_bvalid(qdma_inst_m_axib_bvalid),
    .m_axib_bready(qdma_inst_m_axib_bready),
    .m_axib_arid(qdma_inst_m_axib_arid),
    .m_axib_araddr(qdma_inst_m_axib_araddr),
    .m_axib_arlen(qdma_inst_m_axib_arlen),
    .m_axib_arsize(qdma_inst_m_axib_arsize),
    .m_axib_arburst(qdma_inst_m_axib_arburst),
    .m_axib_arprot(qdma_inst_m_axib_arprot),
    .m_axib_arlock(qdma_inst_m_axib_arlock),
    .m_axib_arcache(qdma_inst_m_axib_arcache),
    .m_axib_arvalid(qdma_inst_m_axib_arvalid),
    .m_axib_arready(qdma_inst_m_axib_arready),
    .m_axib_rid(qdma_inst_m_axib_rid),
    .m_axib_rdata(qdma_inst_m_axib_rdata),
    .m_axib_rresp(qdma_inst_m_axib_rresp),
    .m_axib_rlast(qdma_inst_m_axib_rlast),
    .m_axib_rvalid(qdma_inst_m_axib_rvalid),
    .m_axib_rready(qdma_inst_m_axib_rready),
    .m_axil_awaddr(qdma_inst_m_axil_awaddr),
    .m_axil_awvalid(qdma_inst_m_axil_awvalid),
    .m_axil_awready(qdma_inst_m_axil_awready),
    .m_axil_wdata(qdma_inst_m_axil_wdata),
    .m_axil_wstrb(qdma_inst_m_axil_wstrb),
    .m_axil_wvalid(qdma_inst_m_axil_wvalid),
    .m_axil_wready(qdma_inst_m_axil_wready),
    .m_axil_bresp(qdma_inst_m_axil_bresp),
    .m_axil_bvalid(qdma_inst_m_axil_bvalid),
    .m_axil_bready(qdma_inst_m_axil_bready),
    .m_axil_araddr(qdma_inst_m_axil_araddr),
    .m_axil_arvalid(qdma_inst_m_axil_arvalid),
    .m_axil_arready(qdma_inst_m_axil_arready),
    .m_axil_rdata(qdma_inst_m_axil_rdata),
    .m_axil_rresp(qdma_inst_m_axil_rresp),
    .m_axil_rvalid(qdma_inst_m_axil_rvalid),
    .m_axil_rready(qdma_inst_m_axil_rready),
    .axi_aclk(qdma_inst_axi_aclk),
    .axi_aresetn(qdma_inst_axi_aresetn),
    .soft_reset_n(qdma_inst_soft_reset_n),
    .h2c_byp_in_st_addr(qdma_inst_h2c_byp_in_st_addr),
    .h2c_byp_in_st_len(qdma_inst_h2c_byp_in_st_len),
    .h2c_byp_in_st_eop(qdma_inst_h2c_byp_in_st_eop),
    .h2c_byp_in_st_sop(qdma_inst_h2c_byp_in_st_sop),
    .h2c_byp_in_st_mrkr_req(qdma_inst_h2c_byp_in_st_mrkr_req),
    .h2c_byp_in_st_sdi(qdma_inst_h2c_byp_in_st_sdi),
    .h2c_byp_in_st_qid(qdma_inst_h2c_byp_in_st_qid),
    .h2c_byp_in_st_error(qdma_inst_h2c_byp_in_st_error),
    .h2c_byp_in_st_func(qdma_inst_h2c_byp_in_st_func),
    .h2c_byp_in_st_cidx(qdma_inst_h2c_byp_in_st_cidx),
    .h2c_byp_in_st_port_id(qdma_inst_h2c_byp_in_st_port_id),
    .h2c_byp_in_st_no_dma(qdma_inst_h2c_byp_in_st_no_dma),
    .h2c_byp_in_st_vld(qdma_inst_h2c_byp_in_st_vld),
    .h2c_byp_in_st_rdy(qdma_inst_h2c_byp_in_st_rdy),
    .c2h_byp_in_st_csh_addr(qdma_inst_c2h_byp_in_st_csh_addr),
    .c2h_byp_in_st_csh_qid(qdma_inst_c2h_byp_in_st_csh_qid),
    .c2h_byp_in_st_csh_error(qdma_inst_c2h_byp_in_st_csh_error),
    .c2h_byp_in_st_csh_func(qdma_inst_c2h_byp_in_st_csh_func),
    .c2h_byp_in_st_csh_port_id(qdma_inst_c2h_byp_in_st_csh_port_id),
    .c2h_byp_in_st_csh_pfch_tag(qdma_inst_c2h_byp_in_st_csh_pfch_tag),
    .c2h_byp_in_st_csh_vld(qdma_inst_c2h_byp_in_st_csh_vld),
    .c2h_byp_in_st_csh_rdy(qdma_inst_c2h_byp_in_st_csh_rdy),
    .s_axis_c2h_tdata(qdma_inst_s_axis_c2h_tdata),
    .s_axis_c2h_tcrc(qdma_inst_s_axis_c2h_tcrc),
    .s_axis_c2h_ctrl_marker(qdma_inst_s_axis_c2h_ctrl_marker),
    .s_axis_c2h_ctrl_ecc(qdma_inst_s_axis_c2h_ctrl_ecc),
    .s_axis_c2h_ctrl_len(qdma_inst_s_axis_c2h_ctrl_len),
    .s_axis_c2h_ctrl_port_id(qdma_inst_s_axis_c2h_ctrl_port_id),
    .s_axis_c2h_ctrl_qid(qdma_inst_s_axis_c2h_ctrl_qid),
    .s_axis_c2h_ctrl_has_cmpt(qdma_inst_s_axis_c2h_ctrl_has_cmpt),
    .s_axis_c2h_mty(qdma_inst_s_axis_c2h_mty),
    .s_axis_c2h_tlast(qdma_inst_s_axis_c2h_tlast),
    .s_axis_c2h_tvalid(qdma_inst_s_axis_c2h_tvalid),
    .s_axis_c2h_tready(qdma_inst_s_axis_c2h_tready),
    .m_axis_h2c_tdata(qdma_inst_m_axis_h2c_tdata),
    .m_axis_h2c_tcrc(qdma_inst_m_axis_h2c_tcrc),
    .m_axis_h2c_tuser_qid(qdma_inst_m_axis_h2c_tuser_qid),
    .m_axis_h2c_tuser_port_id(qdma_inst_m_axis_h2c_tuser_port_id),
    .m_axis_h2c_tuser_err(qdma_inst_m_axis_h2c_tuser_err),
    .m_axis_h2c_tuser_mdata(qdma_inst_m_axis_h2c_tuser_mdata),
    .m_axis_h2c_tuser_mty(qdma_inst_m_axis_h2c_tuser_mty),
    .m_axis_h2c_tuser_zero_byte(qdma_inst_m_axis_h2c_tuser_zero_byte),
    .m_axis_h2c_tlast(qdma_inst_m_axis_h2c_tlast),
    .m_axis_h2c_tvalid(qdma_inst_m_axis_h2c_tvalid),
    .m_axis_h2c_tready(qdma_inst_m_axis_h2c_tready),
    .axis_c2h_status_drop(qdma_inst_axis_c2h_status_drop),
    .axis_c2h_status_last(qdma_inst_axis_c2h_status_last),
    .axis_c2h_status_cmp(qdma_inst_axis_c2h_status_cmp),
    .axis_c2h_status_valid(qdma_inst_axis_c2h_status_valid),
    .axis_c2h_status_error(qdma_inst_axis_c2h_status_error),
    .axis_c2h_status_qid(qdma_inst_axis_c2h_status_qid),
    .s_axis_c2h_cmpt_tdata(qdma_inst_s_axis_c2h_cmpt_tdata),
    .s_axis_c2h_cmpt_size(qdma_inst_s_axis_c2h_cmpt_size),
    .s_axis_c2h_cmpt_dpar(qdma_inst_s_axis_c2h_cmpt_dpar),
    .s_axis_c2h_cmpt_tvalid(qdma_inst_s_axis_c2h_cmpt_tvalid),
    .s_axis_c2h_cmpt_tready(qdma_inst_s_axis_c2h_cmpt_tready),
    .s_axis_c2h_cmpt_ctrl_qid(qdma_inst_s_axis_c2h_cmpt_ctrl_qid),
    .s_axis_c2h_cmpt_ctrl_cmpt_type(qdma_inst_s_axis_c2h_cmpt_ctrl_cmpt_type),
    .s_axis_c2h_cmpt_ctrl_wait_pld_pkt_id(qdma_inst_s_axis_c2h_cmpt_ctrl_wait_pld_pkt_id),
    .s_axis_c2h_cmpt_ctrl_no_wrb_marker(qdma_inst_s_axis_c2h_cmpt_ctrl_no_wrb_marker),
    .s_axis_c2h_cmpt_ctrl_port_id(qdma_inst_s_axis_c2h_cmpt_ctrl_port_id),
    .s_axis_c2h_cmpt_ctrl_marker(qdma_inst_s_axis_c2h_cmpt_ctrl_marker),
    .s_axis_c2h_cmpt_ctrl_user_trig(qdma_inst_s_axis_c2h_cmpt_ctrl_user_trig),
    .s_axis_c2h_cmpt_ctrl_col_idx(qdma_inst_s_axis_c2h_cmpt_ctrl_col_idx),
    .s_axis_c2h_cmpt_ctrl_err_idx(qdma_inst_s_axis_c2h_cmpt_ctrl_err_idx),
    .h2c_byp_out_rdy(qdma_inst_h2c_byp_out_rdy),
    .c2h_byp_out_rdy(qdma_inst_c2h_byp_out_rdy),
    .tm_dsc_sts_rdy(qdma_inst_tm_dsc_sts_rdy),
    .dsc_crdt_in_vld(qdma_inst_dsc_crdt_in_vld),
    .dsc_crdt_in_rdy(qdma_inst_dsc_crdt_in_rdy),
    .dsc_crdt_in_dir(qdma_inst_dsc_crdt_in_dir),
    .dsc_crdt_in_fence(qdma_inst_dsc_crdt_in_fence),
    .dsc_crdt_in_qid(qdma_inst_dsc_crdt_in_qid),
    .dsc_crdt_in_crdt(qdma_inst_dsc_crdt_in_crdt),
    .qsts_out_rdy(qdma_inst_qsts_out_rdy),
    .usr_irq_in_vld(qdma_inst_usr_irq_in_vld),
    .usr_irq_in_vec(qdma_inst_usr_irq_in_vec),
    .usr_irq_in_fnc(qdma_inst_usr_irq_in_fnc),
    .usr_irq_out_ack(qdma_inst_usr_irq_out_ack),
    .usr_irq_out_fail(qdma_inst_usr_irq_out_fail)
  );
  assign io_pin_tx_p = qdma_inst_pci_exp_txp; // @[QDMA.scala 139:57]
  assign io_pin_tx_n = qdma_inst_pci_exp_txn; // @[QDMA.scala 138:57]
  assign io_pcie_clk = qdma_inst_axi_aclk; // @[QDMA.scala 143:57]
  assign io_pcie_arstn = qdma_inst_axi_aresetn; // @[QDMA.scala 144:57]
  assign io_h2c_cmd_ready = check_h2c_io_in_ready; // @[QDMA.scala 87:41]
  assign io_h2c_data_valid = fifo_h2c_data_io_out_valid; // @[QDMA.scala 78:33]
  assign io_h2c_data_bits_data = fifo_h2c_data_io_out_bits_data; // @[QDMA.scala 78:33]
  assign io_c2h_cmd_ready = check_c2h_io_in_ready; // @[QDMA.scala 85:41]
  assign io_c2h_data_ready = boundary_split_io_data_in_ready; // @[QDMA.scala 128:41]
  assign io_reg_control_8 = axil2reg_io_reg_control_8; // @[QDMA.scala 111:33]
  assign io_reg_control_9 = axil2reg_io_reg_control_9; // @[QDMA.scala 111:33]
  assign io_reg_control_10 = axil2reg_io_reg_control_10; // @[QDMA.scala 111:33]
  assign io_reg_control_11 = axil2reg_io_reg_control_11; // @[QDMA.scala 111:33]
  assign io_reg_control_12 = axil2reg_io_reg_control_12; // @[QDMA.scala 111:33]
  assign io_reg_control_13 = axil2reg_io_reg_control_13; // @[QDMA.scala 111:33]
  assign io_reg_control_20 = axil2reg_io_reg_control_20; // @[QDMA.scala 111:33]
  assign io_reg_control_50 = axil2reg_io_reg_control_50; // @[QDMA.scala 111:33]
  assign io_reg_control_51 = axil2reg_io_reg_control_51; // @[QDMA.scala 111:33]
  assign io_reg_control_52 = axil2reg_io_reg_control_52; // @[QDMA.scala 111:33]
  assign io_reg_control_53 = axil2reg_io_reg_control_53; // @[QDMA.scala 111:33]
  assign io_reg_control_54 = axil2reg_io_reg_control_54; // @[QDMA.scala 111:33]
  assign io_reg_control_55 = axil2reg_io_reg_control_55; // @[QDMA.scala 111:33]
  assign io_reg_control_56 = axil2reg_io_reg_control_56; // @[QDMA.scala 111:33]
  assign io_reg_control_57 = axil2reg_io_reg_control_57; // @[QDMA.scala 111:33]
  assign io_reg_control_58 = axil2reg_io_reg_control_58; // @[QDMA.scala 111:33]
  assign io_reg_control_59 = axil2reg_io_reg_control_59; // @[QDMA.scala 111:33]
  assign io_reg_control_70 = axil2reg_io_reg_control_70; // @[QDMA.scala 111:33]
  assign io_reg_control_71 = axil2reg_io_reg_control_71; // @[QDMA.scala 111:33]
  assign io_reg_control_72 = axil2reg_io_reg_control_72; // @[QDMA.scala 111:33]
  assign io_reg_control_73 = axil2reg_io_reg_control_73; // @[QDMA.scala 111:33]
  assign io_reg_control_74 = axil2reg_io_reg_control_74; // @[QDMA.scala 111:33]
  assign io_reg_control_75 = axil2reg_io_reg_control_75; // @[QDMA.scala 111:33]
  assign io_reg_control_76 = axil2reg_io_reg_control_76; // @[QDMA.scala 111:33]
  assign io_reg_control_77 = axil2reg_io_reg_control_77; // @[QDMA.scala 111:33]
  assign io_reg_control_78 = axil2reg_io_reg_control_78; // @[QDMA.scala 111:33]
  assign io_reg_control_79 = axil2reg_io_reg_control_79; // @[QDMA.scala 111:33]
  assign io_reg_control_80 = axil2reg_io_reg_control_80; // @[QDMA.scala 111:33]
  assign io_reg_control_91 = axil2reg_io_reg_control_91; // @[QDMA.scala 111:33]
  assign io_reg_control_92 = axil2reg_io_reg_control_92; // @[QDMA.scala 111:33]
  assign io_reg_control_93 = axil2reg_io_reg_control_93; // @[QDMA.scala 111:33]
  assign io_reg_control_94 = axil2reg_io_reg_control_94; // @[QDMA.scala 111:33]
  assign io_axib_aw_valid = qdma_inst_m_axib_awvalid; // @[QDMA.scala 215:65]
  assign io_axib_aw_bits_addr = qdma_inst_m_axib_awaddr; // @[QDMA.scala 208:65]
  assign io_axib_aw_bits_burst = qdma_inst_m_axib_awburst; // @[QDMA.scala 211:65]
  assign io_axib_aw_bits_len = qdma_inst_m_axib_awlen; // @[QDMA.scala 209:65]
  assign io_axib_aw_bits_size = qdma_inst_m_axib_awsize; // @[QDMA.scala 210:65]
  assign io_axib_ar_valid = qdma_inst_m_axib_arvalid; // @[QDMA.scala 237:65]
  assign io_axib_ar_bits_addr = qdma_inst_m_axib_araddr; // @[QDMA.scala 230:65]
  assign io_axib_ar_bits_burst = qdma_inst_m_axib_arburst; // @[QDMA.scala 233:65]
  assign io_axib_ar_bits_len = qdma_inst_m_axib_arlen; // @[QDMA.scala 231:65]
  assign io_axib_ar_bits_size = qdma_inst_m_axib_arsize; // @[QDMA.scala 232:65]
  assign io_axib_w_valid = qdma_inst_m_axib_wvalid; // @[QDMA.scala 221:65]
  assign io_axib_w_bits_data = qdma_inst_m_axib_wdata; // @[QDMA.scala 218:65]
  assign io_axib_w_bits_last = qdma_inst_m_axib_wlast; // @[QDMA.scala 220:65]
  assign io_axib_w_bits_strb = qdma_inst_m_axib_wstrb; // @[QDMA.scala 219:65]
  assign io_axib_r_ready = qdma_inst_m_axib_rready; // @[QDMA.scala 245:65]
  assign io_c2h_status_last = qdma_inst_axis_c2h_status_last; // @[QDMA.scala 188:57]
  assign io_c2h_status_cmp = qdma_inst_axis_c2h_status_cmp; // @[QDMA.scala 189:57]
  assign io_c2h_status_valid = qdma_inst_axis_c2h_status_valid; // @[QDMA.scala 190:57]
  assign io_c2h_status_error = qdma_inst_axis_c2h_status_error; // @[QDMA.scala 191:57]
  assign io_c2h_status_drop = qdma_inst_axis_c2h_status_drop; // @[QDMA.scala 192:57]
  assign io_tlb_miss_count = tlb_io_tlb_miss_count; // @[QDMA.scala 112:41]
  assign perst_n_pad_I = io_pin_sys_rst_n; // @[Buf.scala 18:26]
  assign ibufds_gte4_inst_CEB = 1'h0; // @[QDMA.scala 73:41]
  assign ibufds_gte4_inst_I = io_pin_sys_clk_p; // @[QDMA.scala 72:41]
  assign ibufds_gte4_inst_IB = io_pin_sys_clk_n; // @[QDMA.scala 71:41]
  assign fifo_h2c_data_io_in_clk = io_pcie_clk; // @[XConverter.scala 62:33]
  assign fifo_h2c_data_io_out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign fifo_h2c_data_io_rstn = io_pcie_arstn; // @[XConverter.scala 64:41]
  assign fifo_h2c_data_io_in_valid = qdma_inst_m_axis_h2c_tvalid; // @[QDMA.scala 204:57]
  assign fifo_h2c_data_io_in_bits_data = qdma_inst_m_axis_h2c_tdata; // @[QDMA.scala 195:57]
  assign fifo_h2c_data_io_in_bits_tcrc = qdma_inst_m_axis_h2c_tcrc; // @[QDMA.scala 196:57]
  assign fifo_h2c_data_io_in_bits_tuser_qid = qdma_inst_m_axis_h2c_tuser_qid; // @[QDMA.scala 197:57]
  assign fifo_h2c_data_io_in_bits_tuser_port_id = qdma_inst_m_axis_h2c_tuser_port_id; // @[QDMA.scala 198:49]
  assign fifo_h2c_data_io_in_bits_tuser_err = qdma_inst_m_axis_h2c_tuser_err; // @[QDMA.scala 199:57]
  assign fifo_h2c_data_io_in_bits_tuser_mdata = qdma_inst_m_axis_h2c_tuser_mdata; // @[QDMA.scala 200:57]
  assign fifo_h2c_data_io_in_bits_tuser_mty = qdma_inst_m_axis_h2c_tuser_mty; // @[QDMA.scala 201:57]
  assign fifo_h2c_data_io_in_bits_tuser_zero_byte = qdma_inst_m_axis_h2c_tuser_zero_byte; // @[QDMA.scala 202:49]
  assign fifo_h2c_data_io_in_bits_last = qdma_inst_m_axis_h2c_tlast; // @[QDMA.scala 203:57]
  assign fifo_h2c_data_io_out_ready = io_h2c_data_ready; // @[QDMA.scala 78:33]
  assign fifo_c2h_data_io_in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign fifo_c2h_data_io_out_clk = io_pcie_clk; // @[XConverter.scala 63:33]
  assign fifo_c2h_data_io_rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign fifo_c2h_data_io_in_valid = boundary_split_io_data_out_valid; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_data = boundary_split_io_data_out_bits_data; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_tcrc = boundary_split_io_data_out_bits_tcrc; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_ctrl_marker = boundary_split_io_data_out_bits_ctrl_marker; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_ctrl_ecc = boundary_split_io_data_out_bits_ctrl_ecc; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_ctrl_len = boundary_split_io_data_out_bits_ctrl_len; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_ctrl_port_id = boundary_split_io_data_out_bits_ctrl_port_id; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_ctrl_qid = boundary_split_io_data_out_bits_ctrl_qid; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_ctrl_has_cmpt = boundary_split_io_data_out_bits_ctrl_has_cmpt; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_last = boundary_split_io_data_out_bits_last; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_in_bits_mty = boundary_split_io_data_out_bits_mty; // @[QDMA.scala 130:41]
  assign fifo_c2h_data_io_out_ready = qdma_inst_s_axis_c2h_tready; // @[QDMA.scala 185:57]
  assign fifo_h2c_cmd_io_in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign fifo_h2c_cmd_io_out_clk = io_pcie_clk; // @[XConverter.scala 63:33]
  assign fifo_h2c_cmd_io_rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign fifo_h2c_cmd_io_in_valid = tlb_io_h2c_out_valid; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_addr = tlb_io_h2c_out_bits_addr; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_len = tlb_io_h2c_out_bits_len; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_eop = tlb_io_h2c_out_bits_eop; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_sop = tlb_io_h2c_out_bits_sop; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_mrkr_req = tlb_io_h2c_out_bits_mrkr_req; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_sdi = tlb_io_h2c_out_bits_sdi; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_qid = tlb_io_h2c_out_bits_qid; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_error = tlb_io_h2c_out_bits_error; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_func = tlb_io_h2c_out_bits_func; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_cidx = tlb_io_h2c_out_bits_cidx; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_port_id = tlb_io_h2c_out_bits_port_id; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_in_bits_no_dma = tlb_io_h2c_out_bits_no_dma; // @[QDMA.scala 92:25]
  assign fifo_h2c_cmd_io_out_ready = qdma_inst_h2c_byp_in_st_rdy; // @[QDMA.scala 161:49]
  assign fifo_c2h_cmd_io_in_clk = io_user_clk; // @[XConverter.scala 62:33]
  assign fifo_c2h_cmd_io_out_clk = io_pcie_clk; // @[XConverter.scala 63:33]
  assign fifo_c2h_cmd_io_rstn = io_user_arstn; // @[XConverter.scala 64:41]
  assign fifo_c2h_cmd_io_in_valid = boundary_split_io_cmd_out_valid; // @[QDMA.scala 129:41]
  assign fifo_c2h_cmd_io_in_bits_addr = boundary_split_io_cmd_out_bits_addr; // @[QDMA.scala 129:41]
  assign fifo_c2h_cmd_io_in_bits_qid = boundary_split_io_cmd_out_bits_qid; // @[QDMA.scala 129:41]
  assign fifo_c2h_cmd_io_in_bits_error = boundary_split_io_cmd_out_bits_error; // @[QDMA.scala 129:41]
  assign fifo_c2h_cmd_io_in_bits_func = boundary_split_io_cmd_out_bits_func; // @[QDMA.scala 129:41]
  assign fifo_c2h_cmd_io_in_bits_port_id = boundary_split_io_cmd_out_bits_port_id; // @[QDMA.scala 129:41]
  assign fifo_c2h_cmd_io_in_bits_pfch_tag = boundary_split_io_cmd_out_bits_pfch_tag; // @[QDMA.scala 129:41]
  assign fifo_c2h_cmd_io_in_bits_len = boundary_split_io_cmd_out_bits_len; // @[QDMA.scala 129:41]
  assign fifo_c2h_cmd_io_out_ready = qdma_inst_c2h_byp_in_st_csh_rdy; // @[QDMA.scala 171:57]
  assign check_c2h_clock = io_user_clk;
  assign check_c2h_reset = ~io_user_arstn; // @[QDMA.scala 84:73]
  assign check_c2h_io_in_valid = io_c2h_cmd_valid; // @[QDMA.scala 85:41]
  assign check_c2h_io_in_bits_addr = io_c2h_cmd_bits_addr; // @[QDMA.scala 85:41]
  assign check_c2h_io_in_bits_pfch_tag = io_c2h_cmd_bits_pfch_tag; // @[QDMA.scala 85:41]
  assign check_c2h_io_in_bits_len = io_c2h_cmd_bits_len; // @[QDMA.scala 85:41]
  assign check_c2h_io_out_ready = tlb_io_c2h_in_ready; // @[QDMA.scala 91:25]
  assign check_h2c_clock = io_user_clk;
  assign check_h2c_reset = ~io_user_arstn; // @[QDMA.scala 86:73]
  assign check_h2c_io_in_valid = io_h2c_cmd_valid; // @[QDMA.scala 87:41]
  assign check_h2c_io_in_bits_addr = io_h2c_cmd_bits_addr; // @[QDMA.scala 87:41]
  assign check_h2c_io_in_bits_len = io_h2c_cmd_bits_len; // @[QDMA.scala 87:41]
  assign check_h2c_io_out_ready = tlb_io_h2c_in_ready; // @[QDMA.scala 90:25]
  assign tlb_clock = io_user_clk;
  assign tlb_reset = ~io_user_arstn; // @[QDMA.scala 89:65]
  assign tlb_io_wr_tlb_valid = fifo_wr_tlb_io_out_valid; // @[QDMA.scala 105:41]
  assign tlb_io_wr_tlb_bits_vaddr_high = fifo_wr_tlb_io_out_bits_vaddr_high; // @[QDMA.scala 104:49]
  assign tlb_io_wr_tlb_bits_vaddr_low = fifo_wr_tlb_io_out_bits_vaddr_low; // @[QDMA.scala 104:49]
  assign tlb_io_wr_tlb_bits_paddr_high = fifo_wr_tlb_io_out_bits_paddr_high; // @[QDMA.scala 104:49]
  assign tlb_io_wr_tlb_bits_paddr_low = fifo_wr_tlb_io_out_bits_paddr_low; // @[QDMA.scala 104:49]
  assign tlb_io_wr_tlb_bits_is_base = fifo_wr_tlb_io_out_bits_is_base; // @[QDMA.scala 104:49]
  assign tlb_io_h2c_in_valid = check_h2c_io_out_valid; // @[QDMA.scala 90:25]
  assign tlb_io_h2c_in_bits_addr = check_h2c_io_out_bits_addr; // @[QDMA.scala 90:25]
  assign tlb_io_h2c_in_bits_len = check_h2c_io_out_bits_len; // @[QDMA.scala 90:25]
  assign tlb_io_h2c_in_bits_eop = check_h2c_io_out_bits_eop; // @[QDMA.scala 90:25]
  assign tlb_io_h2c_in_bits_sop = check_h2c_io_out_bits_sop; // @[QDMA.scala 90:25]
  assign tlb_io_c2h_in_valid = check_c2h_io_out_valid; // @[QDMA.scala 91:25]
  assign tlb_io_c2h_in_bits_addr = check_c2h_io_out_bits_addr; // @[QDMA.scala 91:25]
  assign tlb_io_c2h_in_bits_pfch_tag = check_c2h_io_out_bits_pfch_tag; // @[QDMA.scala 91:25]
  assign tlb_io_c2h_in_bits_len = check_c2h_io_out_bits_len; // @[QDMA.scala 91:25]
  assign tlb_io_h2c_out_ready = fifo_h2c_cmd_io_in_ready; // @[QDMA.scala 92:25]
  assign tlb_io_c2h_out_ready = boundary_split_io_cmd_in_ready; // @[QDMA.scala 127:41]
  assign fifo_wr_tlb_io_in_clk = io_pcie_clk; // @[XConverter.scala 62:33]
  assign fifo_wr_tlb_io_out_clk = io_user_clk; // @[XConverter.scala 63:33]
  assign fifo_wr_tlb_io_rstn = io_pcie_arstn; // @[XConverter.scala 64:41]
  assign fifo_wr_tlb_io_in_valid = fifo_wr_tlb_io_in_valid_REG_1; // @[QDMA.scala 102:41]
  assign fifo_wr_tlb_io_in_bits_vaddr_high = io_reg_control_9; // @[QDMA.scala 99:49]
  assign fifo_wr_tlb_io_in_bits_vaddr_low = io_reg_control_8; // @[QDMA.scala 100:49]
  assign fifo_wr_tlb_io_in_bits_paddr_high = io_reg_control_11; // @[QDMA.scala 97:49]
  assign fifo_wr_tlb_io_in_bits_paddr_low = io_reg_control_10; // @[QDMA.scala 98:49]
  assign fifo_wr_tlb_io_in_bits_is_base = io_reg_control_12[0]; // @[QDMA.scala 96:70]
  assign axil2reg_clock = io_pcie_clk;
  assign axil2reg_reset = ~io_pcie_arstn; // @[QDMA.scala 108:54]
  assign axil2reg_io_axi_aw_valid = qdma_inst_m_axil_awvalid; // @[QDMA.scala 249:65]
  assign axil2reg_io_axi_aw_bits_addr = qdma_inst_m_axil_awaddr; // @[QDMA.scala 248:65]
  assign axil2reg_io_axi_ar_valid = qdma_inst_m_axil_arvalid; // @[QDMA.scala 262:65]
  assign axil2reg_io_axi_ar_bits_addr = qdma_inst_m_axil_araddr; // @[QDMA.scala 261:65]
  assign axil2reg_io_axi_w_valid = qdma_inst_m_axil_wvalid; // @[QDMA.scala 254:65]
  assign axil2reg_io_axi_w_bits_data = qdma_inst_m_axil_wdata; // @[QDMA.scala 252:65]
  assign axil2reg_io_axi_r_ready = qdma_inst_m_axil_rready; // @[QDMA.scala 268:65]
  assign axil2reg_io_reg_status_40 = io_reg_status_40; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_51 = io_reg_status_51; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_52 = io_reg_status_52; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_61 = io_reg_status_61; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_71 = io_reg_status_71; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_72 = io_reg_status_72; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_75 = io_reg_status_75; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_76 = io_reg_status_76; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_77 = io_reg_status_77; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_78 = io_reg_status_78; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_79 = io_reg_status_79; // @[QDMA.scala 110:33]
  assign axil2reg_io_reg_status_81 = io_reg_status_81; // @[QDMA.scala 110:33]
  assign boundary_split_clock = io_user_clk;
  assign boundary_split_reset = ~io_user_arstn; // @[QDMA.scala 126:81]
  assign boundary_split_io_data_in_valid = io_c2h_data_valid; // @[QDMA.scala 128:41]
  assign boundary_split_io_data_in_bits_data = io_c2h_data_bits_data; // @[QDMA.scala 128:41]
  assign boundary_split_io_cmd_in_valid = tlb_io_c2h_out_valid; // @[QDMA.scala 127:41]
  assign boundary_split_io_cmd_in_bits_addr = tlb_io_c2h_out_bits_addr; // @[QDMA.scala 127:41]
  assign boundary_split_io_cmd_in_bits_qid = tlb_io_c2h_out_bits_qid; // @[QDMA.scala 127:41]
  assign boundary_split_io_cmd_in_bits_error = tlb_io_c2h_out_bits_error; // @[QDMA.scala 127:41]
  assign boundary_split_io_cmd_in_bits_func = tlb_io_c2h_out_bits_func; // @[QDMA.scala 127:41]
  assign boundary_split_io_cmd_in_bits_port_id = tlb_io_c2h_out_bits_port_id; // @[QDMA.scala 127:41]
  assign boundary_split_io_cmd_in_bits_pfch_tag = tlb_io_c2h_out_bits_pfch_tag; // @[QDMA.scala 127:41]
  assign boundary_split_io_cmd_in_bits_len = tlb_io_c2h_out_bits_len; // @[QDMA.scala 127:41]
  assign boundary_split_io_data_out_ready = fifo_c2h_data_io_in_ready; // @[QDMA.scala 130:41]
  assign boundary_split_io_cmd_out_ready = fifo_c2h_cmd_io_in_ready; // @[QDMA.scala 129:41]
  assign qdma_inst_sys_rst_n = perst_n_pad_O; // @[QDMA.scala 134:57]
  assign qdma_inst_sys_clk = ibufds_gte4_inst_ODIV2; // @[QDMA.scala 135:57]
  assign qdma_inst_sys_clk_gt = ibufds_gte4_inst_O; // @[QDMA.scala 136:57]
  assign qdma_inst_pci_exp_rxn = io_pin_rx_n; // @[QDMA.scala 140:57]
  assign qdma_inst_pci_exp_rxp = io_pin_rx_p; // @[QDMA.scala 141:57]
  assign qdma_inst_m_axib_awready = io_axib_aw_ready; // @[QDMA.scala 216:65]
  assign qdma_inst_m_axib_wready = io_axib_w_ready; // @[QDMA.scala 222:65]
  assign qdma_inst_m_axib_bid = 4'h0; // @[QDMA.scala 224:65]
  assign qdma_inst_m_axib_bresp = 2'h0; // @[QDMA.scala 225:65]
  assign qdma_inst_m_axib_bvalid = io_axib_b_valid; // @[QDMA.scala 226:65]
  assign qdma_inst_m_axib_arready = io_axib_ar_ready; // @[QDMA.scala 238:65]
  assign qdma_inst_m_axib_rid = 4'h0; // @[QDMA.scala 240:65]
  assign qdma_inst_m_axib_rdata = io_axib_r_bits_data; // @[QDMA.scala 241:65]
  assign qdma_inst_m_axib_rresp = 2'h0; // @[QDMA.scala 242:65]
  assign qdma_inst_m_axib_rlast = io_axib_r_bits_last; // @[QDMA.scala 243:65]
  assign qdma_inst_m_axib_rvalid = io_axib_r_valid; // @[QDMA.scala 244:65]
  assign qdma_inst_m_axil_awready = axil2reg_io_axi_aw_ready; // @[QDMA.scala 250:65]
  assign qdma_inst_m_axil_wready = axil2reg_io_axi_w_ready; // @[QDMA.scala 255:65]
  assign qdma_inst_m_axil_bresp = 2'h0; // @[QDMA.scala 257:65]
  assign qdma_inst_m_axil_bvalid = 1'h1; // @[QDMA.scala 258:65]
  assign qdma_inst_m_axil_arready = axil2reg_io_axi_ar_ready; // @[QDMA.scala 263:65]
  assign qdma_inst_m_axil_rdata = axil2reg_io_axi_r_bits_data; // @[QDMA.scala 265:65]
  assign qdma_inst_m_axil_rresp = 2'h0; // @[QDMA.scala 266:65]
  assign qdma_inst_m_axil_rvalid = axil2reg_io_axi_r_valid; // @[QDMA.scala 267:65]
  assign qdma_inst_soft_reset_n = 1'h1; // @[QDMA.scala 145:57]
  assign qdma_inst_h2c_byp_in_st_addr = fifo_h2c_cmd_io_out_bits_addr; // @[QDMA.scala 148:49]
  assign qdma_inst_h2c_byp_in_st_len = fifo_h2c_cmd_io_out_bits_len; // @[QDMA.scala 149:49]
  assign qdma_inst_h2c_byp_in_st_eop = fifo_h2c_cmd_io_out_bits_eop; // @[QDMA.scala 150:49]
  assign qdma_inst_h2c_byp_in_st_sop = fifo_h2c_cmd_io_out_bits_sop; // @[QDMA.scala 151:49]
  assign qdma_inst_h2c_byp_in_st_mrkr_req = fifo_h2c_cmd_io_out_bits_mrkr_req; // @[QDMA.scala 152:49]
  assign qdma_inst_h2c_byp_in_st_sdi = fifo_h2c_cmd_io_out_bits_sdi; // @[QDMA.scala 153:49]
  assign qdma_inst_h2c_byp_in_st_qid = fifo_h2c_cmd_io_out_bits_qid; // @[QDMA.scala 154:49]
  assign qdma_inst_h2c_byp_in_st_error = fifo_h2c_cmd_io_out_bits_error; // @[QDMA.scala 155:49]
  assign qdma_inst_h2c_byp_in_st_func = fifo_h2c_cmd_io_out_bits_func; // @[QDMA.scala 156:49]
  assign qdma_inst_h2c_byp_in_st_cidx = fifo_h2c_cmd_io_out_bits_cidx; // @[QDMA.scala 157:49]
  assign qdma_inst_h2c_byp_in_st_port_id = fifo_h2c_cmd_io_out_bits_port_id; // @[QDMA.scala 158:49]
  assign qdma_inst_h2c_byp_in_st_no_dma = fifo_h2c_cmd_io_out_bits_no_dma; // @[QDMA.scala 159:49]
  assign qdma_inst_h2c_byp_in_st_vld = fifo_h2c_cmd_io_out_valid; // @[QDMA.scala 160:49]
  assign qdma_inst_c2h_byp_in_st_csh_addr = fifo_c2h_cmd_io_out_bits_addr; // @[QDMA.scala 164:57]
  assign qdma_inst_c2h_byp_in_st_csh_qid = fifo_c2h_cmd_io_out_bits_qid; // @[QDMA.scala 165:57]
  assign qdma_inst_c2h_byp_in_st_csh_error = fifo_c2h_cmd_io_out_bits_error; // @[QDMA.scala 166:49]
  assign qdma_inst_c2h_byp_in_st_csh_func = fifo_c2h_cmd_io_out_bits_func; // @[QDMA.scala 167:57]
  assign qdma_inst_c2h_byp_in_st_csh_port_id = fifo_c2h_cmd_io_out_bits_port_id; // @[QDMA.scala 168:49]
  assign qdma_inst_c2h_byp_in_st_csh_pfch_tag = fifo_c2h_cmd_io_out_bits_pfch_tag; // @[QDMA.scala 169:49]
  assign qdma_inst_c2h_byp_in_st_csh_vld = fifo_c2h_cmd_io_out_valid; // @[QDMA.scala 170:57]
  assign qdma_inst_s_axis_c2h_tdata = fifo_c2h_data_io_out_bits_data; // @[QDMA.scala 174:57]
  assign qdma_inst_s_axis_c2h_tcrc = fifo_c2h_data_io_out_bits_tcrc; // @[QDMA.scala 175:57]
  assign qdma_inst_s_axis_c2h_ctrl_marker = fifo_c2h_data_io_out_bits_ctrl_marker; // @[QDMA.scala 176:57]
  assign qdma_inst_s_axis_c2h_ctrl_ecc = fifo_c2h_data_io_out_bits_ctrl_ecc; // @[QDMA.scala 177:57]
  assign qdma_inst_s_axis_c2h_ctrl_len = fifo_c2h_data_io_out_bits_ctrl_len; // @[QDMA.scala 178:57]
  assign qdma_inst_s_axis_c2h_ctrl_port_id = fifo_c2h_data_io_out_bits_ctrl_port_id; // @[QDMA.scala 179:49]
  assign qdma_inst_s_axis_c2h_ctrl_qid = fifo_c2h_data_io_out_bits_ctrl_qid; // @[QDMA.scala 180:57]
  assign qdma_inst_s_axis_c2h_ctrl_has_cmpt = fifo_c2h_data_io_out_bits_ctrl_has_cmpt; // @[QDMA.scala 181:49]
  assign qdma_inst_s_axis_c2h_mty = fifo_c2h_data_io_out_bits_mty; // @[QDMA.scala 182:65]
  assign qdma_inst_s_axis_c2h_tlast = fifo_c2h_data_io_out_bits_last; // @[QDMA.scala 183:57]
  assign qdma_inst_s_axis_c2h_tvalid = fifo_c2h_data_io_out_valid; // @[QDMA.scala 184:57]
  assign qdma_inst_m_axis_h2c_tready = fifo_h2c_data_io_in_ready; // @[QDMA.scala 205:57]
  assign qdma_inst_s_axis_c2h_cmpt_tdata = 512'h0; // @[QDMA.scala 304:81]
  assign qdma_inst_s_axis_c2h_cmpt_size = 2'h0; // @[QDMA.scala 305:81]
  assign qdma_inst_s_axis_c2h_cmpt_dpar = 16'h0; // @[QDMA.scala 306:81]
  assign qdma_inst_s_axis_c2h_cmpt_tvalid = 1'h0; // @[QDMA.scala 307:81]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_qid = 11'h0; // @[QDMA.scala 308:73]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_cmpt_type = 2'h0; // @[QDMA.scala 309:73]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_wait_pld_pkt_id = 16'h0; // @[QDMA.scala 310:65]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_no_wrb_marker = 1'h0; // @[QDMA.scala 312:81]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_port_id = 3'h0; // @[QDMA.scala 314:73]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_marker = 1'h0; // @[QDMA.scala 315:73]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_user_trig = 1'h0; // @[QDMA.scala 316:73]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_col_idx = 3'h0; // @[QDMA.scala 317:73]
  assign qdma_inst_s_axis_c2h_cmpt_ctrl_err_idx = 3'h0; // @[QDMA.scala 318:73]
  assign qdma_inst_h2c_byp_out_rdy = 1'h1; // @[QDMA.scala 320:57]
  assign qdma_inst_c2h_byp_out_rdy = 1'h1; // @[QDMA.scala 321:57]
  assign qdma_inst_tm_dsc_sts_rdy = 1'h1; // @[QDMA.scala 322:65]
  assign qdma_inst_dsc_crdt_in_vld = 1'h0; // @[QDMA.scala 324:65]
  assign qdma_inst_dsc_crdt_in_dir = 1'h0; // @[QDMA.scala 325:65]
  assign qdma_inst_dsc_crdt_in_fence = 1'h0; // @[QDMA.scala 326:65]
  assign qdma_inst_dsc_crdt_in_qid = 11'h0; // @[QDMA.scala 327:65]
  assign qdma_inst_dsc_crdt_in_crdt = 16'h0; // @[QDMA.scala 328:65]
  assign qdma_inst_qsts_out_rdy = 1'h1; // @[QDMA.scala 330:73]
  assign qdma_inst_usr_irq_in_vld = 1'h0; // @[QDMA.scala 332:73]
  assign qdma_inst_usr_irq_in_vec = 11'h0; // @[QDMA.scala 333:73]
  assign qdma_inst_usr_irq_in_fnc = 8'h0; // @[QDMA.scala 334:73]
  always @(posedge io_pcie_clk) begin
    fifo_wr_tlb_io_in_valid_REG <= io_reg_control_13[0]; // @[QDMA.scala 102:126]
    fifo_wr_tlb_io_in_valid_REG_1 <= ~fifo_wr_tlb_io_in_valid_REG & io_reg_control_13[0]; // @[QDMA.scala 102:131]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fifo_wr_tlb_io_in_valid_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  fifo_wr_tlb_io_in_valid_REG_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SV_STREAM_FIFO_5(
  input          io_m_clk,
  input          io_s_clk,
  input          io_reset_n,
  input  [231:0] io_in_data,
  input          io_in_valid,
  output [231:0] io_out_data,
  output         io_out_valid,
  input          io_out_ready
);
  wire [231:0] meta_m_axis_tdata; // @[Meta.scala 30:26]
  wire [28:0] meta_m_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_m_axis_tlast; // @[Meta.scala 30:26]
  wire  meta_m_axis_tvalid; // @[Meta.scala 30:26]
  wire [6:0] meta_rd_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_s_axis_tready; // @[Meta.scala 30:26]
  wire [6:0] meta_wr_data_count_axis; // @[Meta.scala 30:26]
  wire  meta_m_aclk; // @[Meta.scala 30:26]
  wire  meta_m_axis_tready; // @[Meta.scala 30:26]
  wire  meta_s_aclk; // @[Meta.scala 30:26]
  wire  meta_s_aresetn; // @[Meta.scala 30:26]
  wire [231:0] meta_s_axis_tdata; // @[Meta.scala 30:26]
  wire  meta_s_axis_tdest; // @[Meta.scala 30:26]
  wire  meta_s_axis_tid; // @[Meta.scala 30:26]
  wire [28:0] meta_s_axis_tkeep; // @[Meta.scala 30:26]
  wire  meta_s_axis_tlast; // @[Meta.scala 30:26]
  wire [28:0] meta_s_axis_tstrb; // @[Meta.scala 30:26]
  wire  meta_s_axis_tuser; // @[Meta.scala 30:26]
  wire  meta_s_axis_tvalid; // @[Meta.scala 30:26]
  xpm_fifo_axis
    #(.RD_DATA_COUNT_WIDTH(7), .CLOCKING_MODE("common_clock"), .PACKET_FIFO("false"), .USE_ADV_FEATURES("0404"), .TID_WIDTH(1), .TDEST_WIDTH(1), .PROG_EMPTY_THRESH(10), .TUSER_WIDTH(1), .FIFO_DEPTH(64), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(7), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("auto"), .PROG_FULL_THRESH(10), .TDATA_WIDTH(232), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    meta ( // @[Meta.scala 30:26]
    .m_axis_tdata(meta_m_axis_tdata),
    .m_axis_tkeep(meta_m_axis_tkeep),
    .m_axis_tlast(meta_m_axis_tlast),
    .m_axis_tvalid(meta_m_axis_tvalid),
    .rd_data_count_axis(meta_rd_data_count_axis),
    .s_axis_tready(meta_s_axis_tready),
    .wr_data_count_axis(meta_wr_data_count_axis),
    .m_aclk(meta_m_aclk),
    .m_axis_tready(meta_m_axis_tready),
    .s_aclk(meta_s_aclk),
    .s_aresetn(meta_s_aresetn),
    .s_axis_tdata(meta_s_axis_tdata),
    .s_axis_tdest(meta_s_axis_tdest),
    .s_axis_tid(meta_s_axis_tid),
    .s_axis_tkeep(meta_s_axis_tkeep),
    .s_axis_tlast(meta_s_axis_tlast),
    .s_axis_tstrb(meta_s_axis_tstrb),
    .s_axis_tuser(meta_s_axis_tuser),
    .s_axis_tvalid(meta_s_axis_tvalid)
  );
  assign io_out_data = meta_m_axis_tdata; // @[Meta.scala 31:41]
  assign io_out_valid = meta_m_axis_tvalid; // @[Meta.scala 32:41]
  assign meta_m_aclk = io_m_clk; // @[Meta.scala 37:49]
  assign meta_m_axis_tready = io_out_ready; // @[Meta.scala 38:41]
  assign meta_s_aclk = io_s_clk; // @[Meta.scala 39:49]
  assign meta_s_aresetn = io_reset_n; // @[Meta.scala 40:49]
  assign meta_s_axis_tdata = io_in_data; // @[Meta.scala 41:41]
  assign meta_s_axis_tdest = 1'h0; // @[Meta.scala 42:41]
  assign meta_s_axis_tid = 1'h0; // @[Meta.scala 43:49]
  assign meta_s_axis_tkeep = 29'h1fffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tlast = 1'h1; // @[Meta.scala 45:41]
  assign meta_s_axis_tstrb = 29'h1fffffff; // @[Bitwise.scala 72:12]
  assign meta_s_axis_tuser = 1'h0; // @[Meta.scala 47:41]
  assign meta_s_axis_tvalid = io_in_valid; // @[Meta.scala 48:41]
endmodule
module XQueue_2(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_h2c_start_addr,
  input  [33:0] io_in_bits_h2m_start_addr,
  input  [31:0] io_in_bits_h2m_length,
  input  [31:0] io_in_bits_pkt_size,
  input  [63:0] io_in_bits_h2c_cpt_addr,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_h2c_start_addr,
  output [33:0] io_out_bits_h2m_start_addr,
  output [31:0] io_out_bits_h2m_length,
  output [31:0] io_out_bits_pkt_size,
  output [63:0] io_out_bits_h2c_cpt_addr
);
  wire  fifo_io_m_clk; // @[XQueue.scala 67:42]
  wire  fifo_io_s_clk; // @[XQueue.scala 67:42]
  wire  fifo_io_reset_n; // @[XQueue.scala 67:42]
  wire [231:0] fifo_io_in_data; // @[XQueue.scala 67:42]
  wire  fifo_io_in_valid; // @[XQueue.scala 67:42]
  wire [231:0] fifo_io_out_data; // @[XQueue.scala 67:42]
  wire  fifo_io_out_valid; // @[XQueue.scala 67:42]
  wire  fifo_io_out_ready; // @[XQueue.scala 67:42]
  wire [225:0] _fifo_io_in_data_T = {io_in_bits_h2c_start_addr,io_in_bits_h2m_start_addr,io_in_bits_h2m_length,
    io_in_bits_pkt_size,io_in_bits_h2c_cpt_addr}; // @[XQueue.scala 73:71]
  SV_STREAM_FIFO_5 fifo ( // @[XQueue.scala 67:42]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_out_valid = fifo_io_out_valid; // @[XQueue.scala 78:49]
  assign io_out_bits_h2c_start_addr = fifo_io_out_data[225:162]; // @[XQueue.scala 77:85]
  assign io_out_bits_h2m_start_addr = fifo_io_out_data[161:128]; // @[XQueue.scala 77:85]
  assign io_out_bits_h2m_length = fifo_io_out_data[127:96]; // @[XQueue.scala 77:85]
  assign io_out_bits_pkt_size = fifo_io_out_data[95:64]; // @[XQueue.scala 77:85]
  assign io_out_bits_h2c_cpt_addr = fifo_io_out_data[63:0]; // @[XQueue.scala 77:85]
  assign fifo_io_m_clk = clock; // @[XQueue.scala 70:49]
  assign fifo_io_s_clk = clock; // @[XQueue.scala 69:49]
  assign fifo_io_reset_n = ~reset; // @[XQueue.scala 71:52]
  assign fifo_io_in_data = {{6'd0}, _fifo_io_in_data_T}; // @[XQueue.scala 73:71]
  assign fifo_io_in_valid = io_in_valid; // @[XQueue.scala 74:49]
  assign fifo_io_out_ready = io_out_ready; // @[XQueue.scala 79:49]
endmodule
module h2dcmdqueuehead(
  input         clock,
  input         reset,
  output        io_cmd_in_ready,
  input         io_cmd_in_valid,
  input  [63:0] io_cmd_in_bits_h2c_start_addr,
  input  [33:0] io_cmd_in_bits_h2m_start_addr,
  input  [31:0] io_cmd_in_bits_h2m_length,
  input  [31:0] io_cmd_in_bits_pkt_size,
  input  [63:0] io_cmd_in_bits_h2c_cpt_addr,
  input         io_cmd_out_ready,
  output        io_cmd_out_valid,
  output [63:0] io_cmd_out_bits_h2c_start_addr,
  output [33:0] io_cmd_out_bits_h2m_start_addr,
  output [31:0] io_cmd_out_bits_h2m_length,
  output [63:0] io_cmd_out_bits_h2c_cpt_addr,
  output [31:0] io_h2c_length,
  output        io_h2m_complete,
  input         io_h2m_cpt_complete,
  output        io_last,
  output        io_h2m_last,
  output        io_working,
  output        io_continue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg  cmd_in_ready; // @[h2dcmdqueuehead.scala 23:46]
  reg  cmd_out_valid; // @[h2dcmdqueuehead.scala 24:46]
  reg  h2m_complete; // @[h2dcmdqueuehead.scala 25:46]
  reg  working; // @[h2dcmdqueuehead.scala 26:46]
  reg  last; // @[h2dcmdqueuehead.scala 27:46]
  reg  h2m_last; // @[h2dcmdqueuehead.scala 28:46]
  reg  continue_; // @[h2dcmdqueuehead.scala 29:46]
  reg [31:0] length; // @[h2dcmdqueuehead.scala 38:46]
  reg [63:0] h2c_addr; // @[h2dcmdqueuehead.scala 39:46]
  reg [33:0] h2m_addr; // @[h2dcmdqueuehead.scala 40:46]
  reg [33:0] next_addr; // @[h2dcmdqueuehead.scala 43:46]
  reg [33:0] end_addr; // @[h2dcmdqueuehead.scala 44:46]
  reg [63:0] h2c_cpt_addr; // @[h2dcmdqueuehead.scala 45:46]
  reg [31:0] pkt_size; // @[h2dcmdqueuehead.scala 46:46]
  wire  _T = io_cmd_in_ready & io_cmd_in_valid; // @[Decoupled.scala 40:37]
  wire [33:0] _GEN_40 = {{2'd0}, io_cmd_in_bits_h2m_length}; // @[h2dcmdqueuehead.scala 59:70]
  wire [33:0] _end_addr_T_1 = io_cmd_in_bits_h2m_start_addr + _GEN_40; // @[h2dcmdqueuehead.scala 59:70]
  wire [33:0] _GEN_41 = {{2'd0}, io_cmd_in_bits_pkt_size}; // @[h2dcmdqueuehead.scala 65:70]
  wire [33:0] _next_addr_T_1 = io_cmd_in_bits_h2m_start_addr + _GEN_41; // @[h2dcmdqueuehead.scala 65:70]
  wire [31:0] _GEN_0 = io_cmd_in_bits_h2m_length > io_cmd_in_bits_pkt_size ? io_cmd_in_bits_pkt_size :
    io_cmd_in_bits_h2m_length; // @[h2dcmdqueuehead.scala 62:67 h2dcmdqueuehead.scala 63:37 h2dcmdqueuehead.scala 68:37]
  wire [33:0] _GEN_1 = io_cmd_in_bits_h2m_length > io_cmd_in_bits_pkt_size ? _next_addr_T_1 : _end_addr_T_1; // @[h2dcmdqueuehead.scala 62:67 h2dcmdqueuehead.scala 65:37 h2dcmdqueuehead.scala 70:37]
  wire [63:0] _GEN_3 = _T ? io_cmd_in_bits_h2c_start_addr : h2c_addr; // @[h2dcmdqueuehead.scala 55:27 h2dcmdqueuehead.scala 56:37 h2dcmdqueuehead.scala 39:46]
  wire [33:0] _GEN_4 = _T ? io_cmd_in_bits_h2m_start_addr : h2m_addr; // @[h2dcmdqueuehead.scala 55:27 h2dcmdqueuehead.scala 57:37 h2dcmdqueuehead.scala 40:46]
  wire [31:0] _GEN_8 = _T ? _GEN_0 : length; // @[h2dcmdqueuehead.scala 55:27 h2dcmdqueuehead.scala 38:46]
  wire [33:0] _GEN_9 = _T ? _GEN_1 : next_addr; // @[h2dcmdqueuehead.scala 55:27 h2dcmdqueuehead.scala 43:46]
  wire  _GEN_11 = _T ? 1'h0 : cmd_in_ready; // @[h2dcmdqueuehead.scala 55:27 h2dcmdqueuehead.scala 72:37 h2dcmdqueuehead.scala 23:46]
  wire  _GEN_12 = _T | cmd_out_valid; // @[h2dcmdqueuehead.scala 55:27 h2dcmdqueuehead.scala 73:37 h2dcmdqueuehead.scala 24:46]
  wire  _GEN_13 = _T | working; // @[h2dcmdqueuehead.scala 55:27 h2dcmdqueuehead.scala 74:37 h2dcmdqueuehead.scala 26:46]
  wire  _T_2 = io_cmd_out_ready & io_cmd_out_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_43 = {{32'd0}, length}; // @[h2dcmdqueuehead.scala 87:49]
  wire [63:0] _h2c_addr_T_1 = h2c_addr + _GEN_43; // @[h2dcmdqueuehead.scala 87:49]
  wire [33:0] _GEN_44 = {{2'd0}, length}; // @[h2dcmdqueuehead.scala 88:49]
  wire [33:0] _h2m_addr_T_1 = h2m_addr + _GEN_44; // @[h2dcmdqueuehead.scala 88:49]
  wire [33:0] _T_5 = next_addr + _GEN_44; // @[h2dcmdqueuehead.scala 89:29]
  wire [33:0] _length_T_1 = end_addr - next_addr; // @[h2dcmdqueuehead.scala 94:49]
  wire [33:0] _GEN_14 = _T_5 < end_addr ? {{2'd0}, pkt_size} : _length_T_1; // @[h2dcmdqueuehead.scala 89:49 h2dcmdqueuehead.scala 90:37 h2dcmdqueuehead.scala 94:37]
  wire  _GEN_18 = next_addr == end_addr | last; // @[h2dcmdqueuehead.scala 80:38 h2dcmdqueuehead.scala 82:37 h2dcmdqueuehead.scala 27:46]
  wire  _GEN_20 = next_addr == end_addr ? 1'h0 : 1'h1; // @[h2dcmdqueuehead.scala 80:38 h2dcmdqueuehead.scala 84:37 h2dcmdqueuehead.scala 86:37]
  wire [33:0] _GEN_23 = next_addr == end_addr ? {{2'd0}, _GEN_8} : _GEN_14; // @[h2dcmdqueuehead.scala 80:38]
  wire  _GEN_28 = _T_2 ? _GEN_20 : continue_; // @[h2dcmdqueuehead.scala 77:28 h2dcmdqueuehead.scala 29:46]
  wire [33:0] _GEN_31 = _T_2 ? _GEN_23 : {{2'd0}, _GEN_8}; // @[h2dcmdqueuehead.scala 77:28]
  wire  _GEN_33 = continue_ ? 1'h0 : _GEN_28; // @[h2dcmdqueuehead.scala 101:20 h2dcmdqueuehead.scala 102:25]
  wire  _GEN_34 = last & io_cmd_out_ready | h2m_complete; // @[h2dcmdqueuehead.scala 105:35 h2dcmdqueuehead.scala 106:25 h2dcmdqueuehead.scala 25:46]
  wire  _GEN_37 = last & h2m_complete & io_h2m_cpt_complete | _GEN_11; // @[h2dcmdqueuehead.scala 109:53 h2dcmdqueuehead.scala 112:25]
  wire  _GEN_39 = last & h2m_complete & io_h2m_cpt_complete | _GEN_33; // @[h2dcmdqueuehead.scala 109:53 h2dcmdqueuehead.scala 114:25]
  assign io_cmd_in_ready = cmd_in_ready; // @[h2dcmdqueuehead.scala 30:37]
  assign io_cmd_out_valid = cmd_out_valid; // @[h2dcmdqueuehead.scala 31:37]
  assign io_cmd_out_bits_h2c_start_addr = h2c_addr; // @[h2dcmdqueuehead.scala 49:37]
  assign io_cmd_out_bits_h2m_start_addr = h2m_addr; // @[h2dcmdqueuehead.scala 50:37]
  assign io_cmd_out_bits_h2m_length = length; // @[h2dcmdqueuehead.scala 47:37]
  assign io_cmd_out_bits_h2c_cpt_addr = h2c_cpt_addr; // @[h2dcmdqueuehead.scala 52:37]
  assign io_h2c_length = length; // @[h2dcmdqueuehead.scala 48:37]
  assign io_h2m_complete = h2m_complete; // @[h2dcmdqueuehead.scala 32:37]
  assign io_last = last; // @[h2dcmdqueuehead.scala 33:37]
  assign io_h2m_last = h2m_last; // @[h2dcmdqueuehead.scala 34:37]
  assign io_working = working; // @[h2dcmdqueuehead.scala 35:37]
  assign io_continue = continue_; // @[h2dcmdqueuehead.scala 36:37]
  always @(posedge clock) begin
    cmd_in_ready <= reset | _GEN_37; // @[h2dcmdqueuehead.scala 23:46 h2dcmdqueuehead.scala 23:46]
    if (reset) begin // @[h2dcmdqueuehead.scala 24:46]
      cmd_out_valid <= 1'h0; // @[h2dcmdqueuehead.scala 24:46]
    end else if (_T_2) begin // @[h2dcmdqueuehead.scala 77:28]
      if (next_addr == end_addr) begin // @[h2dcmdqueuehead.scala 80:38]
        cmd_out_valid <= 1'h0; // @[h2dcmdqueuehead.scala 81:37]
      end else begin
        cmd_out_valid <= _GEN_12;
      end
    end else begin
      cmd_out_valid <= _GEN_12;
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 25:46]
      h2m_complete <= 1'h0; // @[h2dcmdqueuehead.scala 25:46]
    end else if (last & h2m_complete & io_h2m_cpt_complete) begin // @[h2dcmdqueuehead.scala 109:53]
      h2m_complete <= 1'h0; // @[h2dcmdqueuehead.scala 110:25]
    end else begin
      h2m_complete <= _GEN_34;
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 26:46]
      working <= 1'h0; // @[h2dcmdqueuehead.scala 26:46]
    end else if (last & h2m_complete & io_h2m_cpt_complete) begin // @[h2dcmdqueuehead.scala 109:53]
      working <= 1'h0; // @[h2dcmdqueuehead.scala 113:25]
    end else begin
      working <= _GEN_13;
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 27:46]
      last <= 1'h0; // @[h2dcmdqueuehead.scala 27:46]
    end else if (last & h2m_complete & io_h2m_cpt_complete) begin // @[h2dcmdqueuehead.scala 109:53]
      last <= 1'h0; // @[h2dcmdqueuehead.scala 111:25]
    end else if (_T_2) begin // @[h2dcmdqueuehead.scala 77:28]
      last <= _GEN_18;
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 28:46]
      h2m_last <= 1'h0; // @[h2dcmdqueuehead.scala 28:46]
    end else if (_T_2) begin // @[h2dcmdqueuehead.scala 77:28]
      if (next_addr == end_addr) begin // @[h2dcmdqueuehead.scala 80:38]
        h2m_last <= 1'h0; // @[h2dcmdqueuehead.scala 83:37]
      end else if (_T_5 < end_addr) begin // @[h2dcmdqueuehead.scala 89:49]
        h2m_last <= 1'h0; // @[h2dcmdqueuehead.scala 92:37]
      end else begin
        h2m_last <= 1'h1; // @[h2dcmdqueuehead.scala 96:37]
      end
    end else if (_T) begin // @[h2dcmdqueuehead.scala 55:27]
      if (!(io_cmd_in_bits_h2m_length > io_cmd_in_bits_pkt_size)) begin // @[h2dcmdqueuehead.scala 62:67]
        h2m_last <= 1'h1; // @[h2dcmdqueuehead.scala 67:37]
      end
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 29:46]
      continue_ <= 1'h0; // @[h2dcmdqueuehead.scala 29:46]
    end else begin
      continue_ <= _GEN_39;
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 38:46]
      length <= 32'h0; // @[h2dcmdqueuehead.scala 38:46]
    end else begin
      length <= _GEN_31[31:0];
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 39:46]
      h2c_addr <= 64'h0; // @[h2dcmdqueuehead.scala 39:46]
    end else if (_T_2) begin // @[h2dcmdqueuehead.scala 77:28]
      if (next_addr == end_addr) begin // @[h2dcmdqueuehead.scala 80:38]
        h2c_addr <= _GEN_3;
      end else begin
        h2c_addr <= _h2c_addr_T_1; // @[h2dcmdqueuehead.scala 87:37]
      end
    end else begin
      h2c_addr <= _GEN_3;
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 40:46]
      h2m_addr <= 34'h0; // @[h2dcmdqueuehead.scala 40:46]
    end else if (_T_2) begin // @[h2dcmdqueuehead.scala 77:28]
      if (next_addr == end_addr) begin // @[h2dcmdqueuehead.scala 80:38]
        h2m_addr <= _GEN_4;
      end else begin
        h2m_addr <= _h2m_addr_T_1; // @[h2dcmdqueuehead.scala 88:37]
      end
    end else begin
      h2m_addr <= _GEN_4;
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 43:46]
      next_addr <= 34'h0; // @[h2dcmdqueuehead.scala 43:46]
    end else if (_T_2) begin // @[h2dcmdqueuehead.scala 77:28]
      if (next_addr == end_addr) begin // @[h2dcmdqueuehead.scala 80:38]
        next_addr <= _GEN_9;
      end else if (_T_5 < end_addr) begin // @[h2dcmdqueuehead.scala 89:49]
        next_addr <= _T_5; // @[h2dcmdqueuehead.scala 91:37]
      end else begin
        next_addr <= end_addr; // @[h2dcmdqueuehead.scala 95:37]
      end
    end else begin
      next_addr <= _GEN_9;
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 44:46]
      end_addr <= 34'h0; // @[h2dcmdqueuehead.scala 44:46]
    end else if (_T) begin // @[h2dcmdqueuehead.scala 55:27]
      end_addr <= _end_addr_T_1; // @[h2dcmdqueuehead.scala 59:37]
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 45:46]
      h2c_cpt_addr <= 64'h0; // @[h2dcmdqueuehead.scala 45:46]
    end else if (_T) begin // @[h2dcmdqueuehead.scala 55:27]
      h2c_cpt_addr <= io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueuehead.scala 60:37]
    end
    if (reset) begin // @[h2dcmdqueuehead.scala 46:46]
      pkt_size <= 32'h8000; // @[h2dcmdqueuehead.scala 46:46]
    end else if (_T) begin // @[h2dcmdqueuehead.scala 55:27]
      pkt_size <= io_cmd_in_bits_pkt_size; // @[h2dcmdqueuehead.scala 61:37]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmd_in_ready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cmd_out_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  h2m_complete = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  working = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  last = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  h2m_last = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  continue_ = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  length = _RAND_7[31:0];
  _RAND_8 = {2{`RANDOM}};
  h2c_addr = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  h2m_addr = _RAND_9[33:0];
  _RAND_10 = {2{`RANDOM}};
  next_addr = _RAND_10[33:0];
  _RAND_11 = {2{`RANDOM}};
  end_addr = _RAND_11[33:0];
  _RAND_12 = {2{`RANDOM}};
  h2c_cpt_addr = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  pkt_size = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module h2dcmdqueue(
  input         clock,
  input         reset,
  input         io_cmd_in_valid,
  input  [63:0] io_cmd_in_bits_h2c_start_addr,
  input  [33:0] io_cmd_in_bits_h2m_start_addr,
  input  [31:0] io_cmd_in_bits_h2m_length,
  input  [31:0] io_cmd_in_bits_pkt_size,
  input  [63:0] io_cmd_in_bits_h2c_cpt_addr,
  input  [31:0] io_qin,
  input         io_cmd_out_ready,
  output        io_cmd_out_valid,
  output [63:0] io_cmd_out_bits_h2c_start_addr,
  output [33:0] io_cmd_out_bits_h2m_start_addr,
  output [31:0] io_cmd_out_bits_h2m_length,
  output [63:0] io_cmd_out_bits_h2c_cpt_addr,
  output [31:0] io_h2c_length,
  output        io_h2m_complete,
  input         io_h2m_cpt_complete,
  output        io_last,
  output        io_h2m_last,
  output [31:0] io_counter
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  Q_0_clock; // @[XQueue.scala 35:23]
  wire  Q_0_reset; // @[XQueue.scala 35:23]
  wire  Q_0_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_0_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_0_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_0_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_0_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_0_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_0_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_0_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_0_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_0_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_0_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_0_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_0_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_1_clock; // @[XQueue.scala 35:23]
  wire  Q_1_reset; // @[XQueue.scala 35:23]
  wire  Q_1_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_1_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_1_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_1_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_1_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_1_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_1_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_1_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_1_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_1_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_1_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_1_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_1_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_2_clock; // @[XQueue.scala 35:23]
  wire  Q_2_reset; // @[XQueue.scala 35:23]
  wire  Q_2_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_2_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_2_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_2_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_2_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_2_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_2_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_2_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_2_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_2_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_2_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_2_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_2_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_3_clock; // @[XQueue.scala 35:23]
  wire  Q_3_reset; // @[XQueue.scala 35:23]
  wire  Q_3_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_3_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_3_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_3_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_3_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_3_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_3_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_3_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_3_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_3_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_3_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_3_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_3_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_4_clock; // @[XQueue.scala 35:23]
  wire  Q_4_reset; // @[XQueue.scala 35:23]
  wire  Q_4_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_4_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_4_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_4_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_4_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_4_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_4_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_4_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_4_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_4_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_4_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_4_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_4_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_5_clock; // @[XQueue.scala 35:23]
  wire  Q_5_reset; // @[XQueue.scala 35:23]
  wire  Q_5_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_5_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_5_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_5_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_5_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_5_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_5_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_5_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_5_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_5_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_5_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_5_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_5_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_6_clock; // @[XQueue.scala 35:23]
  wire  Q_6_reset; // @[XQueue.scala 35:23]
  wire  Q_6_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_6_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_6_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_6_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_6_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_6_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_6_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_6_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_6_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_6_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_6_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_6_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_6_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_7_clock; // @[XQueue.scala 35:23]
  wire  Q_7_reset; // @[XQueue.scala 35:23]
  wire  Q_7_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_7_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_7_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_7_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_7_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_7_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_7_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_7_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_7_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_7_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_7_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_7_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_7_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_8_clock; // @[XQueue.scala 35:23]
  wire  Q_8_reset; // @[XQueue.scala 35:23]
  wire  Q_8_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_8_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_8_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_8_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_8_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_8_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_8_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_8_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_8_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_8_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_8_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_8_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_8_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_9_clock; // @[XQueue.scala 35:23]
  wire  Q_9_reset; // @[XQueue.scala 35:23]
  wire  Q_9_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_9_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_9_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_9_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_9_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_9_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_9_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_9_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_9_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_9_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_9_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_9_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_9_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_10_clock; // @[XQueue.scala 35:23]
  wire  Q_10_reset; // @[XQueue.scala 35:23]
  wire  Q_10_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_10_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_10_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_10_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_10_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_10_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_10_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_10_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_10_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_10_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_10_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_10_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_10_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_11_clock; // @[XQueue.scala 35:23]
  wire  Q_11_reset; // @[XQueue.scala 35:23]
  wire  Q_11_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_11_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_11_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_11_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_11_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_11_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_11_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_11_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_11_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_11_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_11_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_11_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_11_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_12_clock; // @[XQueue.scala 35:23]
  wire  Q_12_reset; // @[XQueue.scala 35:23]
  wire  Q_12_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_12_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_12_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_12_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_12_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_12_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_12_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_12_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_12_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_12_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_12_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_12_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_12_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_13_clock; // @[XQueue.scala 35:23]
  wire  Q_13_reset; // @[XQueue.scala 35:23]
  wire  Q_13_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_13_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_13_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_13_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_13_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_13_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_13_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_13_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_13_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_13_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_13_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_13_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_13_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_14_clock; // @[XQueue.scala 35:23]
  wire  Q_14_reset; // @[XQueue.scala 35:23]
  wire  Q_14_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_14_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_14_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_14_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_14_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_14_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_14_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_14_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_14_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_14_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_14_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_14_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_14_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_15_clock; // @[XQueue.scala 35:23]
  wire  Q_15_reset; // @[XQueue.scala 35:23]
  wire  Q_15_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_15_io_in_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_15_io_in_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_15_io_in_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_15_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_15_io_in_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Q_15_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_15_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_15_io_out_bits_h2c_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_15_io_out_bits_h2m_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_15_io_out_bits_h2m_length; // @[XQueue.scala 35:23]
  wire [31:0] Q_15_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire [63:0] Q_15_io_out_bits_h2c_cpt_addr; // @[XQueue.scala 35:23]
  wire  Qh_0_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_0_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_0_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_0_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_0_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_0_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_0_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_0_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_0_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_0_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_0_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_0_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_1_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_1_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_1_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_1_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_1_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_1_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_1_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_1_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_1_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_1_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_1_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_2_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_2_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_2_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_2_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_2_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_2_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_2_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_2_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_2_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_2_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_2_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_3_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_3_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_3_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_3_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_3_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_3_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_3_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_3_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_3_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_3_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_3_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_4_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_4_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_4_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_4_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_4_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_4_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_4_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_4_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_4_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_4_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_4_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_5_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_5_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_5_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_5_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_5_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_5_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_5_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_5_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_5_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_5_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_5_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_6_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_6_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_6_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_6_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_6_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_6_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_6_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_6_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_6_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_6_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_6_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_7_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_7_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_7_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_7_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_7_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_7_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_7_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_7_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_7_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_7_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_7_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_8_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_8_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_8_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_8_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_8_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_8_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_8_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_8_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_8_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_8_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_8_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_9_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_9_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_9_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_9_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_9_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_9_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_9_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_9_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_9_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_9_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_9_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_10_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_10_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_10_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_10_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_10_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_10_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_10_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_10_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_10_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_10_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_10_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_11_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_11_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_11_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_11_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_11_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_11_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_11_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_11_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_11_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_11_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_11_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_12_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_12_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_12_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_12_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_12_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_12_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_12_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_12_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_12_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_12_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_12_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_13_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_13_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_13_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_13_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_13_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_13_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_13_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_13_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_13_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_13_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_13_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_14_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_14_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_14_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_14_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_14_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_14_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_14_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_14_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_14_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_14_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_14_io_continue; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_clock; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_reset; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_cmd_in_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_cmd_in_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_15_io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_15_io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_15_io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_15_io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_15_io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_cmd_out_ready; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_cmd_out_valid; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_15_io_cmd_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [33:0] Qh_15_io_cmd_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_15_io_cmd_out_bits_h2m_length; // @[h2dcmdqueue.scala 27:45]
  wire [63:0] Qh_15_io_cmd_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 27:45]
  wire [31:0] Qh_15_io_h2c_length; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_h2m_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_h2m_cpt_complete; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_h2m_last; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_working; // @[h2dcmdqueue.scala 27:45]
  wire  Qh_15_io_continue; // @[h2dcmdqueue.scala 27:45]
  reg [31:0] counter; // @[h2dcmdqueue.scala 29:26]
  wire  _T = io_cmd_out_ready & io_cmd_out_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[h2dcmdqueue.scala 33:28]
  reg [4:0] out; // @[h2dcmdqueue.scala 36:23]
  reg [4:0] next; // @[h2dcmdqueue.scala 37:23]
  wire  _Qh_0_io_cmd_out_ready_T = out == 5'h0; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_1_io_cmd_out_ready_T = out == 5'h1; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_2_io_cmd_out_ready_T = out == 5'h2; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_3_io_cmd_out_ready_T = out == 5'h3; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_4_io_cmd_out_ready_T = out == 5'h4; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_5_io_cmd_out_ready_T = out == 5'h5; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_6_io_cmd_out_ready_T = out == 5'h6; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_7_io_cmd_out_ready_T = out == 5'h7; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_8_io_cmd_out_ready_T = out == 5'h8; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_9_io_cmd_out_ready_T = out == 5'h9; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_10_io_cmd_out_ready_T = out == 5'ha; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_11_io_cmd_out_ready_T = out == 5'hb; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_12_io_cmd_out_ready_T = out == 5'hc; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_13_io_cmd_out_ready_T = out == 5'hd; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_14_io_cmd_out_ready_T = out == 5'he; // @[h2dcmdqueue.scala 43:64]
  wire  _Qh_15_io_cmd_out_ready_T = out == 5'hf; // @[h2dcmdqueue.scala 43:64]
  wire  _T_1 = ~Qh_0_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_1 = ~Qh_0_io_working & _Qh_0_io_cmd_out_ready_T ? next : out; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17 h2dcmdqueue.scala 36:23]
  wire [4:0] _T_8 = 5'h10 - 5'h1; // @[h2dcmdqueue.scala 55:36]
  wire [4:0] _next_T_1 = next + 5'h1; // @[h2dcmdqueue.scala 58:30]
  wire [4:0] _GEN_2 = next == _T_8 ? 5'h0 : _next_T_1; // @[h2dcmdqueue.scala 55:42 h2dcmdqueue.scala 56:22 h2dcmdqueue.scala 58:22]
  wire [4:0] _GEN_3 = Qh_0_io_continue & _Qh_0_io_cmd_out_ready_T ? next : _GEN_1; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_4 = Qh_0_io_continue & _Qh_0_io_cmd_out_ready_T ? _GEN_2 : next; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 37:23]
  wire [4:0] _GEN_6 = _T_1 & next == 5'h0 ? _GEN_2 : _GEN_4; // @[h2dcmdqueue.scala 61:58]
  wire  _T_16 = ~Qh_1_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_7 = ~Qh_1_io_working & _Qh_1_io_cmd_out_ready_T ? next : _GEN_3; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_9 = Qh_1_io_continue & _Qh_1_io_cmd_out_ready_T ? next : _GEN_7; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_10 = Qh_1_io_continue & _Qh_1_io_cmd_out_ready_T ? _GEN_2 : _GEN_6; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_12 = _T_16 & next == 5'h1 ? _GEN_2 : _GEN_10; // @[h2dcmdqueue.scala 61:58]
  wire  _T_31 = ~Qh_2_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_13 = ~Qh_2_io_working & _Qh_2_io_cmd_out_ready_T ? next : _GEN_9; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_15 = Qh_2_io_continue & _Qh_2_io_cmd_out_ready_T ? next : _GEN_13; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_16 = Qh_2_io_continue & _Qh_2_io_cmd_out_ready_T ? _GEN_2 : _GEN_12; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_18 = _T_31 & next == 5'h2 ? _GEN_2 : _GEN_16; // @[h2dcmdqueue.scala 61:58]
  wire  _T_46 = ~Qh_3_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_19 = ~Qh_3_io_working & _Qh_3_io_cmd_out_ready_T ? next : _GEN_15; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_21 = Qh_3_io_continue & _Qh_3_io_cmd_out_ready_T ? next : _GEN_19; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_22 = Qh_3_io_continue & _Qh_3_io_cmd_out_ready_T ? _GEN_2 : _GEN_18; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_24 = _T_46 & next == 5'h3 ? _GEN_2 : _GEN_22; // @[h2dcmdqueue.scala 61:58]
  wire  _T_61 = ~Qh_4_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_25 = ~Qh_4_io_working & _Qh_4_io_cmd_out_ready_T ? next : _GEN_21; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_27 = Qh_4_io_continue & _Qh_4_io_cmd_out_ready_T ? next : _GEN_25; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_28 = Qh_4_io_continue & _Qh_4_io_cmd_out_ready_T ? _GEN_2 : _GEN_24; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_30 = _T_61 & next == 5'h4 ? _GEN_2 : _GEN_28; // @[h2dcmdqueue.scala 61:58]
  wire  _T_76 = ~Qh_5_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_31 = ~Qh_5_io_working & _Qh_5_io_cmd_out_ready_T ? next : _GEN_27; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_33 = Qh_5_io_continue & _Qh_5_io_cmd_out_ready_T ? next : _GEN_31; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_34 = Qh_5_io_continue & _Qh_5_io_cmd_out_ready_T ? _GEN_2 : _GEN_30; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_36 = _T_76 & next == 5'h5 ? _GEN_2 : _GEN_34; // @[h2dcmdqueue.scala 61:58]
  wire  _T_91 = ~Qh_6_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_37 = ~Qh_6_io_working & _Qh_6_io_cmd_out_ready_T ? next : _GEN_33; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_39 = Qh_6_io_continue & _Qh_6_io_cmd_out_ready_T ? next : _GEN_37; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_40 = Qh_6_io_continue & _Qh_6_io_cmd_out_ready_T ? _GEN_2 : _GEN_36; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_42 = _T_91 & next == 5'h6 ? _GEN_2 : _GEN_40; // @[h2dcmdqueue.scala 61:58]
  wire  _T_106 = ~Qh_7_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_43 = ~Qh_7_io_working & _Qh_7_io_cmd_out_ready_T ? next : _GEN_39; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_45 = Qh_7_io_continue & _Qh_7_io_cmd_out_ready_T ? next : _GEN_43; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_46 = Qh_7_io_continue & _Qh_7_io_cmd_out_ready_T ? _GEN_2 : _GEN_42; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_48 = _T_106 & next == 5'h7 ? _GEN_2 : _GEN_46; // @[h2dcmdqueue.scala 61:58]
  wire  _T_121 = ~Qh_8_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_49 = ~Qh_8_io_working & _Qh_8_io_cmd_out_ready_T ? next : _GEN_45; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_51 = Qh_8_io_continue & _Qh_8_io_cmd_out_ready_T ? next : _GEN_49; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_52 = Qh_8_io_continue & _Qh_8_io_cmd_out_ready_T ? _GEN_2 : _GEN_48; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_54 = _T_121 & next == 5'h8 ? _GEN_2 : _GEN_52; // @[h2dcmdqueue.scala 61:58]
  wire  _T_136 = ~Qh_9_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_55 = ~Qh_9_io_working & _Qh_9_io_cmd_out_ready_T ? next : _GEN_51; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_57 = Qh_9_io_continue & _Qh_9_io_cmd_out_ready_T ? next : _GEN_55; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_58 = Qh_9_io_continue & _Qh_9_io_cmd_out_ready_T ? _GEN_2 : _GEN_54; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_60 = _T_136 & next == 5'h9 ? _GEN_2 : _GEN_58; // @[h2dcmdqueue.scala 61:58]
  wire  _T_151 = ~Qh_10_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_61 = ~Qh_10_io_working & _Qh_10_io_cmd_out_ready_T ? next : _GEN_57; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_63 = Qh_10_io_continue & _Qh_10_io_cmd_out_ready_T ? next : _GEN_61; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_64 = Qh_10_io_continue & _Qh_10_io_cmd_out_ready_T ? _GEN_2 : _GEN_60; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_66 = _T_151 & next == 5'ha ? _GEN_2 : _GEN_64; // @[h2dcmdqueue.scala 61:58]
  wire  _T_166 = ~Qh_11_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_67 = ~Qh_11_io_working & _Qh_11_io_cmd_out_ready_T ? next : _GEN_63; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_69 = Qh_11_io_continue & _Qh_11_io_cmd_out_ready_T ? next : _GEN_67; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_70 = Qh_11_io_continue & _Qh_11_io_cmd_out_ready_T ? _GEN_2 : _GEN_66; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_72 = _T_166 & next == 5'hb ? _GEN_2 : _GEN_70; // @[h2dcmdqueue.scala 61:58]
  wire  _T_181 = ~Qh_12_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_73 = ~Qh_12_io_working & _Qh_12_io_cmd_out_ready_T ? next : _GEN_69; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_75 = Qh_12_io_continue & _Qh_12_io_cmd_out_ready_T ? next : _GEN_73; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_76 = Qh_12_io_continue & _Qh_12_io_cmd_out_ready_T ? _GEN_2 : _GEN_72; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_78 = _T_181 & next == 5'hc ? _GEN_2 : _GEN_76; // @[h2dcmdqueue.scala 61:58]
  wire  _T_196 = ~Qh_13_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_79 = ~Qh_13_io_working & _Qh_13_io_cmd_out_ready_T ? next : _GEN_75; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_81 = Qh_13_io_continue & _Qh_13_io_cmd_out_ready_T ? next : _GEN_79; // @[h2dcmdqueue.scala 53:58 h2dcmdqueue.scala 54:17]
  wire [4:0] _GEN_82 = Qh_13_io_continue & _Qh_13_io_cmd_out_ready_T ? _GEN_2 : _GEN_78; // @[h2dcmdqueue.scala 53:58]
  wire [4:0] _GEN_84 = _T_196 & next == 5'hd ? _GEN_2 : _GEN_82; // @[h2dcmdqueue.scala 61:58]
  wire  _T_211 = ~Qh_14_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [4:0] _GEN_85 = ~Qh_14_io_working & _Qh_14_io_cmd_out_ready_T ? next : _GEN_81; // @[h2dcmdqueue.scala 50:58 h2dcmdqueue.scala 51:17]
  wire [4:0] _GEN_88 = Qh_14_io_continue & _Qh_14_io_cmd_out_ready_T ? _GEN_2 : _GEN_84; // @[h2dcmdqueue.scala 53:58]
  wire  _T_226 = ~Qh_15_io_working; // @[h2dcmdqueue.scala 50:32]
  wire [63:0] _io_cmd_out_bits_T_1_h2c_start_addr = Qh_0_io_cmd_out_bits_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_1_h2m_start_addr = Qh_0_io_cmd_out_bits_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_1_h2m_length = Qh_0_io_cmd_out_bits_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_1_h2c_cpt_addr = Qh_0_io_cmd_out_bits_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_3_h2c_start_addr = 5'h1 == out ? Qh_1_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_1_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_3_h2m_start_addr = 5'h1 == out ? Qh_1_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_1_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_3_h2m_length = 5'h1 == out ? Qh_1_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_1_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_3_h2c_cpt_addr = 5'h1 == out ? Qh_1_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_1_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_5_h2c_start_addr = 5'h2 == out ? Qh_2_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_3_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_5_h2m_start_addr = 5'h2 == out ? Qh_2_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_3_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_5_h2m_length = 5'h2 == out ? Qh_2_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_3_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_5_h2c_cpt_addr = 5'h2 == out ? Qh_2_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_3_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_7_h2c_start_addr = 5'h3 == out ? Qh_3_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_5_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_7_h2m_start_addr = 5'h3 == out ? Qh_3_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_5_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_7_h2m_length = 5'h3 == out ? Qh_3_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_5_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_7_h2c_cpt_addr = 5'h3 == out ? Qh_3_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_5_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_9_h2c_start_addr = 5'h4 == out ? Qh_4_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_7_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_9_h2m_start_addr = 5'h4 == out ? Qh_4_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_7_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_9_h2m_length = 5'h4 == out ? Qh_4_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_7_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_9_h2c_cpt_addr = 5'h4 == out ? Qh_4_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_7_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_11_h2c_start_addr = 5'h5 == out ? Qh_5_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_9_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_11_h2m_start_addr = 5'h5 == out ? Qh_5_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_9_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_11_h2m_length = 5'h5 == out ? Qh_5_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_9_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_11_h2c_cpt_addr = 5'h5 == out ? Qh_5_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_9_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_13_h2c_start_addr = 5'h6 == out ? Qh_6_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_11_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_13_h2m_start_addr = 5'h6 == out ? Qh_6_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_11_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_13_h2m_length = 5'h6 == out ? Qh_6_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_11_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_13_h2c_cpt_addr = 5'h6 == out ? Qh_6_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_11_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_15_h2c_start_addr = 5'h7 == out ? Qh_7_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_13_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_15_h2m_start_addr = 5'h7 == out ? Qh_7_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_13_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_15_h2m_length = 5'h7 == out ? Qh_7_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_13_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_15_h2c_cpt_addr = 5'h7 == out ? Qh_7_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_13_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_17_h2c_start_addr = 5'h8 == out ? Qh_8_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_15_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_17_h2m_start_addr = 5'h8 == out ? Qh_8_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_15_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_17_h2m_length = 5'h8 == out ? Qh_8_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_15_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_17_h2c_cpt_addr = 5'h8 == out ? Qh_8_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_15_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_19_h2c_start_addr = 5'h9 == out ? Qh_9_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_17_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_19_h2m_start_addr = 5'h9 == out ? Qh_9_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_17_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_19_h2m_length = 5'h9 == out ? Qh_9_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_17_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_19_h2c_cpt_addr = 5'h9 == out ? Qh_9_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_17_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_21_h2c_start_addr = 5'ha == out ? Qh_10_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_19_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_21_h2m_start_addr = 5'ha == out ? Qh_10_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_19_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_21_h2m_length = 5'ha == out ? Qh_10_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_19_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_21_h2c_cpt_addr = 5'ha == out ? Qh_10_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_19_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_23_h2c_start_addr = 5'hb == out ? Qh_11_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_21_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_23_h2m_start_addr = 5'hb == out ? Qh_11_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_21_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_23_h2m_length = 5'hb == out ? Qh_11_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_21_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_23_h2c_cpt_addr = 5'hb == out ? Qh_11_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_21_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_25_h2c_start_addr = 5'hc == out ? Qh_12_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_23_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_25_h2m_start_addr = 5'hc == out ? Qh_12_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_23_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_25_h2m_length = 5'hc == out ? Qh_12_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_23_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_25_h2c_cpt_addr = 5'hc == out ? Qh_12_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_23_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_27_h2c_start_addr = 5'hd == out ? Qh_13_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_25_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_27_h2m_start_addr = 5'hd == out ? Qh_13_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_25_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_27_h2m_length = 5'hd == out ? Qh_13_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_25_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_27_h2c_cpt_addr = 5'hd == out ? Qh_13_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_25_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_29_h2c_start_addr = 5'he == out ? Qh_14_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_27_h2c_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_29_h2m_start_addr = 5'he == out ? Qh_14_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_27_h2m_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_29_h2m_length = 5'he == out ? Qh_14_io_cmd_out_bits_h2m_length :
    _io_cmd_out_bits_T_27_h2m_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_29_h2c_cpt_addr = 5'he == out ? Qh_14_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_27_h2c_cpt_addr; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_3 = 5'h1 == out ? Qh_1_io_cmd_out_valid : Qh_0_io_cmd_out_valid; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_5 = 5'h2 == out ? Qh_2_io_cmd_out_valid : _io_cmd_out_valid_T_3; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_7 = 5'h3 == out ? Qh_3_io_cmd_out_valid : _io_cmd_out_valid_T_5; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_9 = 5'h4 == out ? Qh_4_io_cmd_out_valid : _io_cmd_out_valid_T_7; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_11 = 5'h5 == out ? Qh_5_io_cmd_out_valid : _io_cmd_out_valid_T_9; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_13 = 5'h6 == out ? Qh_6_io_cmd_out_valid : _io_cmd_out_valid_T_11; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_15 = 5'h7 == out ? Qh_7_io_cmd_out_valid : _io_cmd_out_valid_T_13; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_17 = 5'h8 == out ? Qh_8_io_cmd_out_valid : _io_cmd_out_valid_T_15; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_19 = 5'h9 == out ? Qh_9_io_cmd_out_valid : _io_cmd_out_valid_T_17; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_21 = 5'ha == out ? Qh_10_io_cmd_out_valid : _io_cmd_out_valid_T_19; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_23 = 5'hb == out ? Qh_11_io_cmd_out_valid : _io_cmd_out_valid_T_21; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_25 = 5'hc == out ? Qh_12_io_cmd_out_valid : _io_cmd_out_valid_T_23; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_27 = 5'hd == out ? Qh_13_io_cmd_out_valid : _io_cmd_out_valid_T_25; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_29 = 5'he == out ? Qh_14_io_cmd_out_valid : _io_cmd_out_valid_T_27; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_1 = Qh_0_io_h2c_length; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_3 = 5'h1 == out ? Qh_1_io_h2c_length : _io_h2c_length_T_1; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_5 = 5'h2 == out ? Qh_2_io_h2c_length : _io_h2c_length_T_3; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_7 = 5'h3 == out ? Qh_3_io_h2c_length : _io_h2c_length_T_5; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_9 = 5'h4 == out ? Qh_4_io_h2c_length : _io_h2c_length_T_7; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_11 = 5'h5 == out ? Qh_5_io_h2c_length : _io_h2c_length_T_9; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_13 = 5'h6 == out ? Qh_6_io_h2c_length : _io_h2c_length_T_11; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_15 = 5'h7 == out ? Qh_7_io_h2c_length : _io_h2c_length_T_13; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_17 = 5'h8 == out ? Qh_8_io_h2c_length : _io_h2c_length_T_15; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_19 = 5'h9 == out ? Qh_9_io_h2c_length : _io_h2c_length_T_17; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_21 = 5'ha == out ? Qh_10_io_h2c_length : _io_h2c_length_T_19; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_23 = 5'hb == out ? Qh_11_io_h2c_length : _io_h2c_length_T_21; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_25 = 5'hc == out ? Qh_12_io_h2c_length : _io_h2c_length_T_23; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_27 = 5'hd == out ? Qh_13_io_h2c_length : _io_h2c_length_T_25; // @[Mux.scala 80:57]
  wire [31:0] _io_h2c_length_T_29 = 5'he == out ? Qh_14_io_h2c_length : _io_h2c_length_T_27; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_3 = 5'h1 == out ? Qh_1_io_h2m_complete : Qh_0_io_h2m_complete; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_5 = 5'h2 == out ? Qh_2_io_h2m_complete : _io_h2m_complete_T_3; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_7 = 5'h3 == out ? Qh_3_io_h2m_complete : _io_h2m_complete_T_5; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_9 = 5'h4 == out ? Qh_4_io_h2m_complete : _io_h2m_complete_T_7; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_11 = 5'h5 == out ? Qh_5_io_h2m_complete : _io_h2m_complete_T_9; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_13 = 5'h6 == out ? Qh_6_io_h2m_complete : _io_h2m_complete_T_11; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_15 = 5'h7 == out ? Qh_7_io_h2m_complete : _io_h2m_complete_T_13; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_17 = 5'h8 == out ? Qh_8_io_h2m_complete : _io_h2m_complete_T_15; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_19 = 5'h9 == out ? Qh_9_io_h2m_complete : _io_h2m_complete_T_17; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_21 = 5'ha == out ? Qh_10_io_h2m_complete : _io_h2m_complete_T_19; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_23 = 5'hb == out ? Qh_11_io_h2m_complete : _io_h2m_complete_T_21; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_25 = 5'hc == out ? Qh_12_io_h2m_complete : _io_h2m_complete_T_23; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_27 = 5'hd == out ? Qh_13_io_h2m_complete : _io_h2m_complete_T_25; // @[Mux.scala 80:57]
  wire  _io_h2m_complete_T_29 = 5'he == out ? Qh_14_io_h2m_complete : _io_h2m_complete_T_27; // @[Mux.scala 80:57]
  wire  _io_last_T_3 = 5'h1 == out ? Qh_1_io_last : Qh_0_io_last; // @[Mux.scala 80:57]
  wire  _io_last_T_5 = 5'h2 == out ? Qh_2_io_last : _io_last_T_3; // @[Mux.scala 80:57]
  wire  _io_last_T_7 = 5'h3 == out ? Qh_3_io_last : _io_last_T_5; // @[Mux.scala 80:57]
  wire  _io_last_T_9 = 5'h4 == out ? Qh_4_io_last : _io_last_T_7; // @[Mux.scala 80:57]
  wire  _io_last_T_11 = 5'h5 == out ? Qh_5_io_last : _io_last_T_9; // @[Mux.scala 80:57]
  wire  _io_last_T_13 = 5'h6 == out ? Qh_6_io_last : _io_last_T_11; // @[Mux.scala 80:57]
  wire  _io_last_T_15 = 5'h7 == out ? Qh_7_io_last : _io_last_T_13; // @[Mux.scala 80:57]
  wire  _io_last_T_17 = 5'h8 == out ? Qh_8_io_last : _io_last_T_15; // @[Mux.scala 80:57]
  wire  _io_last_T_19 = 5'h9 == out ? Qh_9_io_last : _io_last_T_17; // @[Mux.scala 80:57]
  wire  _io_last_T_21 = 5'ha == out ? Qh_10_io_last : _io_last_T_19; // @[Mux.scala 80:57]
  wire  _io_last_T_23 = 5'hb == out ? Qh_11_io_last : _io_last_T_21; // @[Mux.scala 80:57]
  wire  _io_last_T_25 = 5'hc == out ? Qh_12_io_last : _io_last_T_23; // @[Mux.scala 80:57]
  wire  _io_last_T_27 = 5'hd == out ? Qh_13_io_last : _io_last_T_25; // @[Mux.scala 80:57]
  wire  _io_last_T_29 = 5'he == out ? Qh_14_io_last : _io_last_T_27; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_3 = 5'h1 == out ? Qh_1_io_h2m_last : Qh_0_io_h2m_last; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_5 = 5'h2 == out ? Qh_2_io_h2m_last : _io_h2m_last_T_3; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_7 = 5'h3 == out ? Qh_3_io_h2m_last : _io_h2m_last_T_5; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_9 = 5'h4 == out ? Qh_4_io_h2m_last : _io_h2m_last_T_7; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_11 = 5'h5 == out ? Qh_5_io_h2m_last : _io_h2m_last_T_9; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_13 = 5'h6 == out ? Qh_6_io_h2m_last : _io_h2m_last_T_11; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_15 = 5'h7 == out ? Qh_7_io_h2m_last : _io_h2m_last_T_13; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_17 = 5'h8 == out ? Qh_8_io_h2m_last : _io_h2m_last_T_15; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_19 = 5'h9 == out ? Qh_9_io_h2m_last : _io_h2m_last_T_17; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_21 = 5'ha == out ? Qh_10_io_h2m_last : _io_h2m_last_T_19; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_23 = 5'hb == out ? Qh_11_io_h2m_last : _io_h2m_last_T_21; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_25 = 5'hc == out ? Qh_12_io_h2m_last : _io_h2m_last_T_23; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_27 = 5'hd == out ? Qh_13_io_h2m_last : _io_h2m_last_T_25; // @[Mux.scala 80:57]
  wire  _io_h2m_last_T_29 = 5'he == out ? Qh_14_io_h2m_last : _io_h2m_last_T_27; // @[Mux.scala 80:57]
  XQueue_2 Q_0 ( // @[XQueue.scala 35:23]
    .clock(Q_0_clock),
    .reset(Q_0_reset),
    .io_in_valid(Q_0_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_0_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_0_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_0_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_0_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_0_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_0_io_out_ready),
    .io_out_valid(Q_0_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_0_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_0_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_0_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_0_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_0_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_1 ( // @[XQueue.scala 35:23]
    .clock(Q_1_clock),
    .reset(Q_1_reset),
    .io_in_valid(Q_1_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_1_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_1_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_1_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_1_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_1_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_1_io_out_ready),
    .io_out_valid(Q_1_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_1_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_1_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_1_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_1_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_1_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_2 ( // @[XQueue.scala 35:23]
    .clock(Q_2_clock),
    .reset(Q_2_reset),
    .io_in_valid(Q_2_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_2_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_2_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_2_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_2_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_2_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_2_io_out_ready),
    .io_out_valid(Q_2_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_2_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_2_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_2_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_2_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_2_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_3 ( // @[XQueue.scala 35:23]
    .clock(Q_3_clock),
    .reset(Q_3_reset),
    .io_in_valid(Q_3_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_3_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_3_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_3_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_3_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_3_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_3_io_out_ready),
    .io_out_valid(Q_3_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_3_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_3_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_3_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_3_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_3_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_4 ( // @[XQueue.scala 35:23]
    .clock(Q_4_clock),
    .reset(Q_4_reset),
    .io_in_valid(Q_4_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_4_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_4_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_4_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_4_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_4_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_4_io_out_ready),
    .io_out_valid(Q_4_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_4_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_4_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_4_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_4_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_4_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_5 ( // @[XQueue.scala 35:23]
    .clock(Q_5_clock),
    .reset(Q_5_reset),
    .io_in_valid(Q_5_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_5_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_5_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_5_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_5_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_5_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_5_io_out_ready),
    .io_out_valid(Q_5_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_5_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_5_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_5_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_5_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_5_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_6 ( // @[XQueue.scala 35:23]
    .clock(Q_6_clock),
    .reset(Q_6_reset),
    .io_in_valid(Q_6_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_6_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_6_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_6_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_6_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_6_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_6_io_out_ready),
    .io_out_valid(Q_6_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_6_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_6_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_6_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_6_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_6_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_7 ( // @[XQueue.scala 35:23]
    .clock(Q_7_clock),
    .reset(Q_7_reset),
    .io_in_valid(Q_7_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_7_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_7_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_7_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_7_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_7_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_7_io_out_ready),
    .io_out_valid(Q_7_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_7_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_7_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_7_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_7_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_7_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_8 ( // @[XQueue.scala 35:23]
    .clock(Q_8_clock),
    .reset(Q_8_reset),
    .io_in_valid(Q_8_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_8_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_8_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_8_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_8_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_8_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_8_io_out_ready),
    .io_out_valid(Q_8_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_8_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_8_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_8_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_8_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_8_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_9 ( // @[XQueue.scala 35:23]
    .clock(Q_9_clock),
    .reset(Q_9_reset),
    .io_in_valid(Q_9_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_9_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_9_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_9_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_9_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_9_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_9_io_out_ready),
    .io_out_valid(Q_9_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_9_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_9_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_9_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_9_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_9_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_10 ( // @[XQueue.scala 35:23]
    .clock(Q_10_clock),
    .reset(Q_10_reset),
    .io_in_valid(Q_10_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_10_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_10_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_10_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_10_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_10_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_10_io_out_ready),
    .io_out_valid(Q_10_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_10_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_10_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_10_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_10_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_10_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_11 ( // @[XQueue.scala 35:23]
    .clock(Q_11_clock),
    .reset(Q_11_reset),
    .io_in_valid(Q_11_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_11_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_11_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_11_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_11_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_11_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_11_io_out_ready),
    .io_out_valid(Q_11_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_11_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_11_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_11_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_11_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_11_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_12 ( // @[XQueue.scala 35:23]
    .clock(Q_12_clock),
    .reset(Q_12_reset),
    .io_in_valid(Q_12_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_12_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_12_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_12_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_12_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_12_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_12_io_out_ready),
    .io_out_valid(Q_12_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_12_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_12_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_12_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_12_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_12_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_13 ( // @[XQueue.scala 35:23]
    .clock(Q_13_clock),
    .reset(Q_13_reset),
    .io_in_valid(Q_13_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_13_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_13_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_13_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_13_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_13_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_13_io_out_ready),
    .io_out_valid(Q_13_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_13_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_13_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_13_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_13_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_13_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_14 ( // @[XQueue.scala 35:23]
    .clock(Q_14_clock),
    .reset(Q_14_reset),
    .io_in_valid(Q_14_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_14_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_14_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_14_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_14_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_14_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_14_io_out_ready),
    .io_out_valid(Q_14_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_14_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_14_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_14_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_14_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_14_io_out_bits_h2c_cpt_addr)
  );
  XQueue_2 Q_15 ( // @[XQueue.scala 35:23]
    .clock(Q_15_clock),
    .reset(Q_15_reset),
    .io_in_valid(Q_15_io_in_valid),
    .io_in_bits_h2c_start_addr(Q_15_io_in_bits_h2c_start_addr),
    .io_in_bits_h2m_start_addr(Q_15_io_in_bits_h2m_start_addr),
    .io_in_bits_h2m_length(Q_15_io_in_bits_h2m_length),
    .io_in_bits_pkt_size(Q_15_io_in_bits_pkt_size),
    .io_in_bits_h2c_cpt_addr(Q_15_io_in_bits_h2c_cpt_addr),
    .io_out_ready(Q_15_io_out_ready),
    .io_out_valid(Q_15_io_out_valid),
    .io_out_bits_h2c_start_addr(Q_15_io_out_bits_h2c_start_addr),
    .io_out_bits_h2m_start_addr(Q_15_io_out_bits_h2m_start_addr),
    .io_out_bits_h2m_length(Q_15_io_out_bits_h2m_length),
    .io_out_bits_pkt_size(Q_15_io_out_bits_pkt_size),
    .io_out_bits_h2c_cpt_addr(Q_15_io_out_bits_h2c_cpt_addr)
  );
  h2dcmdqueuehead Qh_0 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_0_clock),
    .reset(Qh_0_reset),
    .io_cmd_in_ready(Qh_0_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_0_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_0_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_0_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_0_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_0_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_0_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_0_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_0_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_0_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_0_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_0_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_0_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_0_io_h2c_length),
    .io_h2m_complete(Qh_0_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_0_io_h2m_cpt_complete),
    .io_last(Qh_0_io_last),
    .io_h2m_last(Qh_0_io_h2m_last),
    .io_working(Qh_0_io_working),
    .io_continue(Qh_0_io_continue)
  );
  h2dcmdqueuehead Qh_1 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_1_clock),
    .reset(Qh_1_reset),
    .io_cmd_in_ready(Qh_1_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_1_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_1_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_1_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_1_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_1_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_1_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_1_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_1_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_1_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_1_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_1_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_1_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_1_io_h2c_length),
    .io_h2m_complete(Qh_1_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_1_io_h2m_cpt_complete),
    .io_last(Qh_1_io_last),
    .io_h2m_last(Qh_1_io_h2m_last),
    .io_working(Qh_1_io_working),
    .io_continue(Qh_1_io_continue)
  );
  h2dcmdqueuehead Qh_2 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_2_clock),
    .reset(Qh_2_reset),
    .io_cmd_in_ready(Qh_2_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_2_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_2_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_2_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_2_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_2_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_2_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_2_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_2_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_2_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_2_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_2_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_2_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_2_io_h2c_length),
    .io_h2m_complete(Qh_2_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_2_io_h2m_cpt_complete),
    .io_last(Qh_2_io_last),
    .io_h2m_last(Qh_2_io_h2m_last),
    .io_working(Qh_2_io_working),
    .io_continue(Qh_2_io_continue)
  );
  h2dcmdqueuehead Qh_3 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_3_clock),
    .reset(Qh_3_reset),
    .io_cmd_in_ready(Qh_3_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_3_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_3_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_3_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_3_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_3_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_3_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_3_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_3_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_3_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_3_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_3_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_3_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_3_io_h2c_length),
    .io_h2m_complete(Qh_3_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_3_io_h2m_cpt_complete),
    .io_last(Qh_3_io_last),
    .io_h2m_last(Qh_3_io_h2m_last),
    .io_working(Qh_3_io_working),
    .io_continue(Qh_3_io_continue)
  );
  h2dcmdqueuehead Qh_4 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_4_clock),
    .reset(Qh_4_reset),
    .io_cmd_in_ready(Qh_4_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_4_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_4_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_4_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_4_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_4_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_4_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_4_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_4_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_4_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_4_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_4_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_4_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_4_io_h2c_length),
    .io_h2m_complete(Qh_4_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_4_io_h2m_cpt_complete),
    .io_last(Qh_4_io_last),
    .io_h2m_last(Qh_4_io_h2m_last),
    .io_working(Qh_4_io_working),
    .io_continue(Qh_4_io_continue)
  );
  h2dcmdqueuehead Qh_5 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_5_clock),
    .reset(Qh_5_reset),
    .io_cmd_in_ready(Qh_5_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_5_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_5_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_5_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_5_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_5_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_5_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_5_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_5_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_5_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_5_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_5_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_5_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_5_io_h2c_length),
    .io_h2m_complete(Qh_5_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_5_io_h2m_cpt_complete),
    .io_last(Qh_5_io_last),
    .io_h2m_last(Qh_5_io_h2m_last),
    .io_working(Qh_5_io_working),
    .io_continue(Qh_5_io_continue)
  );
  h2dcmdqueuehead Qh_6 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_6_clock),
    .reset(Qh_6_reset),
    .io_cmd_in_ready(Qh_6_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_6_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_6_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_6_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_6_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_6_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_6_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_6_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_6_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_6_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_6_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_6_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_6_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_6_io_h2c_length),
    .io_h2m_complete(Qh_6_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_6_io_h2m_cpt_complete),
    .io_last(Qh_6_io_last),
    .io_h2m_last(Qh_6_io_h2m_last),
    .io_working(Qh_6_io_working),
    .io_continue(Qh_6_io_continue)
  );
  h2dcmdqueuehead Qh_7 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_7_clock),
    .reset(Qh_7_reset),
    .io_cmd_in_ready(Qh_7_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_7_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_7_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_7_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_7_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_7_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_7_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_7_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_7_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_7_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_7_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_7_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_7_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_7_io_h2c_length),
    .io_h2m_complete(Qh_7_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_7_io_h2m_cpt_complete),
    .io_last(Qh_7_io_last),
    .io_h2m_last(Qh_7_io_h2m_last),
    .io_working(Qh_7_io_working),
    .io_continue(Qh_7_io_continue)
  );
  h2dcmdqueuehead Qh_8 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_8_clock),
    .reset(Qh_8_reset),
    .io_cmd_in_ready(Qh_8_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_8_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_8_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_8_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_8_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_8_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_8_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_8_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_8_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_8_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_8_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_8_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_8_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_8_io_h2c_length),
    .io_h2m_complete(Qh_8_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_8_io_h2m_cpt_complete),
    .io_last(Qh_8_io_last),
    .io_h2m_last(Qh_8_io_h2m_last),
    .io_working(Qh_8_io_working),
    .io_continue(Qh_8_io_continue)
  );
  h2dcmdqueuehead Qh_9 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_9_clock),
    .reset(Qh_9_reset),
    .io_cmd_in_ready(Qh_9_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_9_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_9_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_9_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_9_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_9_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_9_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_9_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_9_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_9_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_9_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_9_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_9_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_9_io_h2c_length),
    .io_h2m_complete(Qh_9_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_9_io_h2m_cpt_complete),
    .io_last(Qh_9_io_last),
    .io_h2m_last(Qh_9_io_h2m_last),
    .io_working(Qh_9_io_working),
    .io_continue(Qh_9_io_continue)
  );
  h2dcmdqueuehead Qh_10 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_10_clock),
    .reset(Qh_10_reset),
    .io_cmd_in_ready(Qh_10_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_10_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_10_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_10_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_10_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_10_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_10_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_10_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_10_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_10_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_10_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_10_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_10_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_10_io_h2c_length),
    .io_h2m_complete(Qh_10_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_10_io_h2m_cpt_complete),
    .io_last(Qh_10_io_last),
    .io_h2m_last(Qh_10_io_h2m_last),
    .io_working(Qh_10_io_working),
    .io_continue(Qh_10_io_continue)
  );
  h2dcmdqueuehead Qh_11 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_11_clock),
    .reset(Qh_11_reset),
    .io_cmd_in_ready(Qh_11_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_11_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_11_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_11_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_11_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_11_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_11_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_11_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_11_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_11_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_11_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_11_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_11_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_11_io_h2c_length),
    .io_h2m_complete(Qh_11_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_11_io_h2m_cpt_complete),
    .io_last(Qh_11_io_last),
    .io_h2m_last(Qh_11_io_h2m_last),
    .io_working(Qh_11_io_working),
    .io_continue(Qh_11_io_continue)
  );
  h2dcmdqueuehead Qh_12 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_12_clock),
    .reset(Qh_12_reset),
    .io_cmd_in_ready(Qh_12_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_12_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_12_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_12_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_12_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_12_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_12_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_12_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_12_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_12_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_12_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_12_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_12_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_12_io_h2c_length),
    .io_h2m_complete(Qh_12_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_12_io_h2m_cpt_complete),
    .io_last(Qh_12_io_last),
    .io_h2m_last(Qh_12_io_h2m_last),
    .io_working(Qh_12_io_working),
    .io_continue(Qh_12_io_continue)
  );
  h2dcmdqueuehead Qh_13 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_13_clock),
    .reset(Qh_13_reset),
    .io_cmd_in_ready(Qh_13_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_13_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_13_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_13_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_13_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_13_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_13_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_13_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_13_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_13_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_13_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_13_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_13_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_13_io_h2c_length),
    .io_h2m_complete(Qh_13_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_13_io_h2m_cpt_complete),
    .io_last(Qh_13_io_last),
    .io_h2m_last(Qh_13_io_h2m_last),
    .io_working(Qh_13_io_working),
    .io_continue(Qh_13_io_continue)
  );
  h2dcmdqueuehead Qh_14 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_14_clock),
    .reset(Qh_14_reset),
    .io_cmd_in_ready(Qh_14_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_14_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_14_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_14_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_14_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_14_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_14_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_14_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_14_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_14_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_14_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_14_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_14_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_14_io_h2c_length),
    .io_h2m_complete(Qh_14_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_14_io_h2m_cpt_complete),
    .io_last(Qh_14_io_last),
    .io_h2m_last(Qh_14_io_h2m_last),
    .io_working(Qh_14_io_working),
    .io_continue(Qh_14_io_continue)
  );
  h2dcmdqueuehead Qh_15 ( // @[h2dcmdqueue.scala 27:45]
    .clock(Qh_15_clock),
    .reset(Qh_15_reset),
    .io_cmd_in_ready(Qh_15_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_15_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(Qh_15_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(Qh_15_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(Qh_15_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(Qh_15_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(Qh_15_io_cmd_in_bits_h2c_cpt_addr),
    .io_cmd_out_ready(Qh_15_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_15_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(Qh_15_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(Qh_15_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(Qh_15_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(Qh_15_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(Qh_15_io_h2c_length),
    .io_h2m_complete(Qh_15_io_h2m_complete),
    .io_h2m_cpt_complete(Qh_15_io_h2m_cpt_complete),
    .io_last(Qh_15_io_last),
    .io_h2m_last(Qh_15_io_h2m_last),
    .io_working(Qh_15_io_working),
    .io_continue(Qh_15_io_continue)
  );
  assign io_cmd_out_valid = 5'hf == out ? Qh_15_io_cmd_out_valid : _io_cmd_out_valid_T_29; // @[Mux.scala 80:57]
  assign io_cmd_out_bits_h2c_start_addr = 5'hf == out ? Qh_15_io_cmd_out_bits_h2c_start_addr :
    _io_cmd_out_bits_T_29_h2c_start_addr; // @[Mux.scala 80:57]
  assign io_cmd_out_bits_h2m_start_addr = 5'hf == out ? Qh_15_io_cmd_out_bits_h2m_start_addr :
    _io_cmd_out_bits_T_29_h2m_start_addr; // @[Mux.scala 80:57]
  assign io_cmd_out_bits_h2m_length = 5'hf == out ? Qh_15_io_cmd_out_bits_h2m_length : _io_cmd_out_bits_T_29_h2m_length; // @[Mux.scala 80:57]
  assign io_cmd_out_bits_h2c_cpt_addr = 5'hf == out ? Qh_15_io_cmd_out_bits_h2c_cpt_addr :
    _io_cmd_out_bits_T_29_h2c_cpt_addr; // @[Mux.scala 80:57]
  assign io_h2c_length = 5'hf == out ? Qh_15_io_h2c_length : _io_h2c_length_T_29; // @[Mux.scala 80:57]
  assign io_h2m_complete = 5'hf == out ? Qh_15_io_h2m_complete : _io_h2m_complete_T_29; // @[Mux.scala 80:57]
  assign io_last = 5'hf == out ? Qh_15_io_last : _io_last_T_29; // @[Mux.scala 80:57]
  assign io_h2m_last = 5'hf == out ? Qh_15_io_h2m_last : _io_h2m_last_T_29; // @[Mux.scala 80:57]
  assign io_counter = counter; // @[h2dcmdqueue.scala 30:16]
  assign Q_0_clock = clock;
  assign Q_0_reset = reset;
  assign Q_0_io_in_valid = io_cmd_in_valid & io_qin[0]; // @[h2dcmdqueue.scala 40:56]
  assign Q_0_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_0_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_0_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_0_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_0_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_0_io_out_ready = Qh_0_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_1_clock = clock;
  assign Q_1_reset = reset;
  assign Q_1_io_in_valid = io_cmd_in_valid & io_qin[1]; // @[h2dcmdqueue.scala 40:56]
  assign Q_1_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_1_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_1_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_1_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_1_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_1_io_out_ready = Qh_1_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_2_clock = clock;
  assign Q_2_reset = reset;
  assign Q_2_io_in_valid = io_cmd_in_valid & io_qin[2]; // @[h2dcmdqueue.scala 40:56]
  assign Q_2_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_2_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_2_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_2_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_2_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_2_io_out_ready = Qh_2_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_3_clock = clock;
  assign Q_3_reset = reset;
  assign Q_3_io_in_valid = io_cmd_in_valid & io_qin[3]; // @[h2dcmdqueue.scala 40:56]
  assign Q_3_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_3_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_3_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_3_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_3_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_3_io_out_ready = Qh_3_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_4_clock = clock;
  assign Q_4_reset = reset;
  assign Q_4_io_in_valid = io_cmd_in_valid & io_qin[4]; // @[h2dcmdqueue.scala 40:56]
  assign Q_4_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_4_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_4_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_4_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_4_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_4_io_out_ready = Qh_4_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_5_clock = clock;
  assign Q_5_reset = reset;
  assign Q_5_io_in_valid = io_cmd_in_valid & io_qin[5]; // @[h2dcmdqueue.scala 40:56]
  assign Q_5_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_5_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_5_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_5_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_5_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_5_io_out_ready = Qh_5_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_6_clock = clock;
  assign Q_6_reset = reset;
  assign Q_6_io_in_valid = io_cmd_in_valid & io_qin[6]; // @[h2dcmdqueue.scala 40:56]
  assign Q_6_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_6_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_6_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_6_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_6_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_6_io_out_ready = Qh_6_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_7_clock = clock;
  assign Q_7_reset = reset;
  assign Q_7_io_in_valid = io_cmd_in_valid & io_qin[7]; // @[h2dcmdqueue.scala 40:56]
  assign Q_7_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_7_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_7_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_7_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_7_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_7_io_out_ready = Qh_7_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_8_clock = clock;
  assign Q_8_reset = reset;
  assign Q_8_io_in_valid = io_cmd_in_valid & io_qin[8]; // @[h2dcmdqueue.scala 40:56]
  assign Q_8_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_8_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_8_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_8_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_8_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_8_io_out_ready = Qh_8_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_9_clock = clock;
  assign Q_9_reset = reset;
  assign Q_9_io_in_valid = io_cmd_in_valid & io_qin[9]; // @[h2dcmdqueue.scala 40:56]
  assign Q_9_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_9_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_9_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_9_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_9_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_9_io_out_ready = Qh_9_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_10_clock = clock;
  assign Q_10_reset = reset;
  assign Q_10_io_in_valid = io_cmd_in_valid & io_qin[10]; // @[h2dcmdqueue.scala 40:56]
  assign Q_10_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_10_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_10_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_10_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_10_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_10_io_out_ready = Qh_10_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_11_clock = clock;
  assign Q_11_reset = reset;
  assign Q_11_io_in_valid = io_cmd_in_valid & io_qin[11]; // @[h2dcmdqueue.scala 40:56]
  assign Q_11_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_11_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_11_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_11_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_11_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_11_io_out_ready = Qh_11_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_12_clock = clock;
  assign Q_12_reset = reset;
  assign Q_12_io_in_valid = io_cmd_in_valid & io_qin[12]; // @[h2dcmdqueue.scala 40:56]
  assign Q_12_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_12_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_12_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_12_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_12_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_12_io_out_ready = Qh_12_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_13_clock = clock;
  assign Q_13_reset = reset;
  assign Q_13_io_in_valid = io_cmd_in_valid & io_qin[13]; // @[h2dcmdqueue.scala 40:56]
  assign Q_13_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_13_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_13_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_13_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_13_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_13_io_out_ready = Qh_13_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_14_clock = clock;
  assign Q_14_reset = reset;
  assign Q_14_io_in_valid = io_cmd_in_valid & io_qin[14]; // @[h2dcmdqueue.scala 40:56]
  assign Q_14_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_14_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_14_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_14_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_14_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_14_io_out_ready = Qh_14_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Q_15_clock = clock;
  assign Q_15_reset = reset;
  assign Q_15_io_in_valid = io_cmd_in_valid & io_qin[15]; // @[h2dcmdqueue.scala 40:56]
  assign Q_15_io_in_bits_h2c_start_addr = io_cmd_in_bits_h2c_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_15_io_in_bits_h2m_start_addr = io_cmd_in_bits_h2m_start_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_15_io_in_bits_h2m_length = io_cmd_in_bits_h2m_length; // @[h2dcmdqueue.scala 41:37]
  assign Q_15_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[h2dcmdqueue.scala 41:37]
  assign Q_15_io_in_bits_h2c_cpt_addr = io_cmd_in_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 41:37]
  assign Q_15_io_out_ready = Qh_15_io_cmd_in_ready; // @[h2dcmdqueue.scala 42:37]
  assign Qh_0_clock = clock;
  assign Qh_0_reset = reset;
  assign Qh_0_io_cmd_in_valid = Q_0_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_0_io_cmd_in_bits_h2c_start_addr = Q_0_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_0_io_cmd_in_bits_h2m_start_addr = Q_0_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_0_io_cmd_in_bits_h2m_length = Q_0_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_0_io_cmd_in_bits_pkt_size = Q_0_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_0_io_cmd_in_bits_h2c_cpt_addr = Q_0_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_0_io_cmd_out_ready = io_cmd_out_ready & out == 5'h0; // @[h2dcmdqueue.scala 43:57]
  assign Qh_0_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_0_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_1_clock = clock;
  assign Qh_1_reset = reset;
  assign Qh_1_io_cmd_in_valid = Q_1_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_1_io_cmd_in_bits_h2c_start_addr = Q_1_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_1_io_cmd_in_bits_h2m_start_addr = Q_1_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_1_io_cmd_in_bits_h2m_length = Q_1_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_1_io_cmd_in_bits_pkt_size = Q_1_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_1_io_cmd_in_bits_h2c_cpt_addr = Q_1_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_1_io_cmd_out_ready = io_cmd_out_ready & out == 5'h1; // @[h2dcmdqueue.scala 43:57]
  assign Qh_1_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_1_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_2_clock = clock;
  assign Qh_2_reset = reset;
  assign Qh_2_io_cmd_in_valid = Q_2_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_2_io_cmd_in_bits_h2c_start_addr = Q_2_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_2_io_cmd_in_bits_h2m_start_addr = Q_2_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_2_io_cmd_in_bits_h2m_length = Q_2_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_2_io_cmd_in_bits_pkt_size = Q_2_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_2_io_cmd_in_bits_h2c_cpt_addr = Q_2_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_2_io_cmd_out_ready = io_cmd_out_ready & out == 5'h2; // @[h2dcmdqueue.scala 43:57]
  assign Qh_2_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_2_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_3_clock = clock;
  assign Qh_3_reset = reset;
  assign Qh_3_io_cmd_in_valid = Q_3_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_3_io_cmd_in_bits_h2c_start_addr = Q_3_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_3_io_cmd_in_bits_h2m_start_addr = Q_3_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_3_io_cmd_in_bits_h2m_length = Q_3_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_3_io_cmd_in_bits_pkt_size = Q_3_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_3_io_cmd_in_bits_h2c_cpt_addr = Q_3_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_3_io_cmd_out_ready = io_cmd_out_ready & out == 5'h3; // @[h2dcmdqueue.scala 43:57]
  assign Qh_3_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_3_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_4_clock = clock;
  assign Qh_4_reset = reset;
  assign Qh_4_io_cmd_in_valid = Q_4_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_4_io_cmd_in_bits_h2c_start_addr = Q_4_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_4_io_cmd_in_bits_h2m_start_addr = Q_4_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_4_io_cmd_in_bits_h2m_length = Q_4_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_4_io_cmd_in_bits_pkt_size = Q_4_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_4_io_cmd_in_bits_h2c_cpt_addr = Q_4_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_4_io_cmd_out_ready = io_cmd_out_ready & out == 5'h4; // @[h2dcmdqueue.scala 43:57]
  assign Qh_4_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_4_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_5_clock = clock;
  assign Qh_5_reset = reset;
  assign Qh_5_io_cmd_in_valid = Q_5_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_5_io_cmd_in_bits_h2c_start_addr = Q_5_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_5_io_cmd_in_bits_h2m_start_addr = Q_5_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_5_io_cmd_in_bits_h2m_length = Q_5_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_5_io_cmd_in_bits_pkt_size = Q_5_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_5_io_cmd_in_bits_h2c_cpt_addr = Q_5_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_5_io_cmd_out_ready = io_cmd_out_ready & out == 5'h5; // @[h2dcmdqueue.scala 43:57]
  assign Qh_5_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_5_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_6_clock = clock;
  assign Qh_6_reset = reset;
  assign Qh_6_io_cmd_in_valid = Q_6_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_6_io_cmd_in_bits_h2c_start_addr = Q_6_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_6_io_cmd_in_bits_h2m_start_addr = Q_6_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_6_io_cmd_in_bits_h2m_length = Q_6_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_6_io_cmd_in_bits_pkt_size = Q_6_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_6_io_cmd_in_bits_h2c_cpt_addr = Q_6_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_6_io_cmd_out_ready = io_cmd_out_ready & out == 5'h6; // @[h2dcmdqueue.scala 43:57]
  assign Qh_6_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_6_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_7_clock = clock;
  assign Qh_7_reset = reset;
  assign Qh_7_io_cmd_in_valid = Q_7_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_7_io_cmd_in_bits_h2c_start_addr = Q_7_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_7_io_cmd_in_bits_h2m_start_addr = Q_7_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_7_io_cmd_in_bits_h2m_length = Q_7_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_7_io_cmd_in_bits_pkt_size = Q_7_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_7_io_cmd_in_bits_h2c_cpt_addr = Q_7_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_7_io_cmd_out_ready = io_cmd_out_ready & out == 5'h7; // @[h2dcmdqueue.scala 43:57]
  assign Qh_7_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_7_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_8_clock = clock;
  assign Qh_8_reset = reset;
  assign Qh_8_io_cmd_in_valid = Q_8_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_8_io_cmd_in_bits_h2c_start_addr = Q_8_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_8_io_cmd_in_bits_h2m_start_addr = Q_8_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_8_io_cmd_in_bits_h2m_length = Q_8_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_8_io_cmd_in_bits_pkt_size = Q_8_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_8_io_cmd_in_bits_h2c_cpt_addr = Q_8_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_8_io_cmd_out_ready = io_cmd_out_ready & out == 5'h8; // @[h2dcmdqueue.scala 43:57]
  assign Qh_8_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_8_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_9_clock = clock;
  assign Qh_9_reset = reset;
  assign Qh_9_io_cmd_in_valid = Q_9_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_9_io_cmd_in_bits_h2c_start_addr = Q_9_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_9_io_cmd_in_bits_h2m_start_addr = Q_9_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_9_io_cmd_in_bits_h2m_length = Q_9_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_9_io_cmd_in_bits_pkt_size = Q_9_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_9_io_cmd_in_bits_h2c_cpt_addr = Q_9_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_9_io_cmd_out_ready = io_cmd_out_ready & out == 5'h9; // @[h2dcmdqueue.scala 43:57]
  assign Qh_9_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_9_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_10_clock = clock;
  assign Qh_10_reset = reset;
  assign Qh_10_io_cmd_in_valid = Q_10_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_10_io_cmd_in_bits_h2c_start_addr = Q_10_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_10_io_cmd_in_bits_h2m_start_addr = Q_10_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_10_io_cmd_in_bits_h2m_length = Q_10_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_10_io_cmd_in_bits_pkt_size = Q_10_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_10_io_cmd_in_bits_h2c_cpt_addr = Q_10_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_10_io_cmd_out_ready = io_cmd_out_ready & out == 5'ha; // @[h2dcmdqueue.scala 43:57]
  assign Qh_10_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_10_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_11_clock = clock;
  assign Qh_11_reset = reset;
  assign Qh_11_io_cmd_in_valid = Q_11_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_11_io_cmd_in_bits_h2c_start_addr = Q_11_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_11_io_cmd_in_bits_h2m_start_addr = Q_11_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_11_io_cmd_in_bits_h2m_length = Q_11_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_11_io_cmd_in_bits_pkt_size = Q_11_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_11_io_cmd_in_bits_h2c_cpt_addr = Q_11_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_11_io_cmd_out_ready = io_cmd_out_ready & out == 5'hb; // @[h2dcmdqueue.scala 43:57]
  assign Qh_11_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_11_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_12_clock = clock;
  assign Qh_12_reset = reset;
  assign Qh_12_io_cmd_in_valid = Q_12_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_12_io_cmd_in_bits_h2c_start_addr = Q_12_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_12_io_cmd_in_bits_h2m_start_addr = Q_12_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_12_io_cmd_in_bits_h2m_length = Q_12_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_12_io_cmd_in_bits_pkt_size = Q_12_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_12_io_cmd_in_bits_h2c_cpt_addr = Q_12_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_12_io_cmd_out_ready = io_cmd_out_ready & out == 5'hc; // @[h2dcmdqueue.scala 43:57]
  assign Qh_12_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_12_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_13_clock = clock;
  assign Qh_13_reset = reset;
  assign Qh_13_io_cmd_in_valid = Q_13_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_13_io_cmd_in_bits_h2c_start_addr = Q_13_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_13_io_cmd_in_bits_h2m_start_addr = Q_13_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_13_io_cmd_in_bits_h2m_length = Q_13_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_13_io_cmd_in_bits_pkt_size = Q_13_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_13_io_cmd_in_bits_h2c_cpt_addr = Q_13_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_13_io_cmd_out_ready = io_cmd_out_ready & out == 5'hd; // @[h2dcmdqueue.scala 43:57]
  assign Qh_13_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_13_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_14_clock = clock;
  assign Qh_14_reset = reset;
  assign Qh_14_io_cmd_in_valid = Q_14_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_14_io_cmd_in_bits_h2c_start_addr = Q_14_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_14_io_cmd_in_bits_h2m_start_addr = Q_14_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_14_io_cmd_in_bits_h2m_length = Q_14_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_14_io_cmd_in_bits_pkt_size = Q_14_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_14_io_cmd_in_bits_h2c_cpt_addr = Q_14_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_14_io_cmd_out_ready = io_cmd_out_ready & out == 5'he; // @[h2dcmdqueue.scala 43:57]
  assign Qh_14_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_14_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  assign Qh_15_clock = clock;
  assign Qh_15_reset = reset;
  assign Qh_15_io_cmd_in_valid = Q_15_io_out_valid; // @[h2dcmdqueue.scala 42:37]
  assign Qh_15_io_cmd_in_bits_h2c_start_addr = Q_15_io_out_bits_h2c_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_15_io_cmd_in_bits_h2m_start_addr = Q_15_io_out_bits_h2m_start_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_15_io_cmd_in_bits_h2m_length = Q_15_io_out_bits_h2m_length; // @[h2dcmdqueue.scala 42:37]
  assign Qh_15_io_cmd_in_bits_pkt_size = Q_15_io_out_bits_pkt_size; // @[h2dcmdqueue.scala 42:37]
  assign Qh_15_io_cmd_in_bits_h2c_cpt_addr = Q_15_io_out_bits_h2c_cpt_addr; // @[h2dcmdqueue.scala 42:37]
  assign Qh_15_io_cmd_out_ready = io_cmd_out_ready & out == 5'hf; // @[h2dcmdqueue.scala 43:57]
  assign Qh_15_io_h2m_cpt_complete = io_h2m_cpt_complete & _Qh_15_io_cmd_out_ready_T; // @[h2dcmdqueue.scala 44:60]
  always @(posedge clock) begin
    if (reset) begin // @[h2dcmdqueue.scala 29:26]
      counter <= 32'h0; // @[h2dcmdqueue.scala 29:26]
    end else if (_T) begin // @[h2dcmdqueue.scala 32:5]
      counter <= _counter_T_1; // @[h2dcmdqueue.scala 33:17]
    end
    if (reset) begin // @[h2dcmdqueue.scala 36:23]
      out <= 5'h0; // @[h2dcmdqueue.scala 36:23]
    end else if (Qh_15_io_continue & _Qh_15_io_cmd_out_ready_T) begin // @[h2dcmdqueue.scala 53:58]
      out <= next; // @[h2dcmdqueue.scala 54:17]
    end else if (~Qh_15_io_working & _Qh_15_io_cmd_out_ready_T) begin // @[h2dcmdqueue.scala 50:58]
      out <= next; // @[h2dcmdqueue.scala 51:17]
    end else if (Qh_14_io_continue & _Qh_14_io_cmd_out_ready_T) begin // @[h2dcmdqueue.scala 53:58]
      out <= next; // @[h2dcmdqueue.scala 54:17]
    end else begin
      out <= _GEN_85;
    end
    if (reset) begin // @[h2dcmdqueue.scala 37:23]
      next <= 5'h0; // @[h2dcmdqueue.scala 37:23]
    end else if (_T_226 & next == 5'hf) begin // @[h2dcmdqueue.scala 61:58]
      next <= _GEN_2;
    end else if (Qh_15_io_continue & _Qh_15_io_cmd_out_ready_T) begin // @[h2dcmdqueue.scala 53:58]
      next <= _GEN_2;
    end else if (_T_211 & next == 5'he) begin // @[h2dcmdqueue.scala 61:58]
      next <= _GEN_2;
    end else begin
      next <= _GEN_88;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  out = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  next = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module H2C(
  input         clock,
  input         reset,
  input  [63:0] io_start_addr,
  input  [31:0] io_length,
  input         io_start,
  input         io_h2c_cmd_ready,
  output        io_h2c_cmd_valid,
  output [63:0] io_h2c_cmd_bits_addr,
  output [31:0] io_h2c_cmd_bits_len,
  output        io_complete,
  output [31:0] io_count_time,
  output [31:0] io_send_cmd_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] addr; // @[H2C.scala 23:50]
  reg [31:0] length; // @[H2C.scala 24:50]
  reg  valid_cmd; // @[H2C.scala 25:42]
  reg [31:0] count_time; // @[H2C.scala 28:42]
  reg [31:0] send_cmd_count; // @[H2C.scala 29:42]
  reg  complete; // @[H2C.scala 32:42]
  reg [3:0] hold; // @[H2C.scala 34:50]
  reg [1:0] state_cmd; // @[H2C.scala 52:42]
  wire  _T = 2'h0 == state_cmd; // @[Conditional.scala 37:30]
  wire  _GEN_1 = io_start ? 1'h0 : complete; // @[H2C.scala 56:39 H2C.scala 58:65 H2C.scala 32:42]
  wire  _T_1 = 2'h1 == state_cmd; // @[Conditional.scala 37:30]
  wire [31:0] _count_time_T_1 = count_time + 32'h1; // @[H2C.scala 67:79]
  wire  _T_2 = io_h2c_cmd_ready & io_h2c_cmd_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = 2'h2 == state_cmd; // @[Conditional.scala 37:30]
  wire [3:0] _hold_T_1 = hold - 4'h1; // @[H2C.scala 76:38]
  wire  _GEN_10 = hold == 4'h0 | complete; // @[H2C.scala 77:44 H2C.scala 78:65 H2C.scala 32:42]
  wire [1:0] _GEN_11 = hold == 4'h0 ? 2'h0 : state_cmd; // @[H2C.scala 77:44 H2C.scala 79:65 H2C.scala 52:42]
  wire  _GEN_13 = _T_3 ? _GEN_10 : complete; // @[Conditional.scala 39:67 H2C.scala 32:42]
  wire  _GEN_19 = _T_1 ? complete : _GEN_13; // @[Conditional.scala 39:67 H2C.scala 32:42]
  wire  _GEN_21 = _T ? _GEN_1 : _GEN_19; // @[Conditional.scala 40:58]
  wire [31:0] _send_cmd_count_T_1 = send_cmd_count + 32'h1; // @[H2C.scala 85:51]
  assign io_h2c_cmd_valid = valid_cmd; // @[H2C.scala 44:33]
  assign io_h2c_cmd_bits_addr = addr; // @[H2C.scala 43:33]
  assign io_h2c_cmd_bits_len = length; // @[H2C.scala 41:33]
  assign io_complete = complete; // @[H2C.scala 88:33]
  assign io_count_time = count_time; // @[H2C.scala 89:33]
  assign io_send_cmd_count = send_cmd_count; // @[H2C.scala 90:33]
  always @(posedge clock) begin
    if (reset) begin // @[H2C.scala 23:50]
      addr <= 64'h0; // @[H2C.scala 23:50]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2C.scala 56:39]
        addr <= io_start_addr; // @[H2C.scala 59:65]
      end
    end
    if (reset) begin // @[H2C.scala 24:50]
      length <= 32'h0; // @[H2C.scala 24:50]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2C.scala 56:39]
        length <= io_length; // @[H2C.scala 60:65]
      end
    end
    if (reset) begin // @[H2C.scala 25:42]
      valid_cmd <= 1'h0; // @[H2C.scala 25:42]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[H2C.scala 69:48]
          valid_cmd <= 1'h0; // @[H2C.scala 71:65]
        end else begin
          valid_cmd <= 1'h1; // @[H2C.scala 68:65]
        end
      end
    end
    if (reset) begin // @[H2C.scala 28:42]
      count_time <= 32'h0; // @[H2C.scala 28:42]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2C.scala 56:39]
        count_time <= 32'h0; // @[H2C.scala 62:65]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      count_time <= _count_time_T_1; // @[H2C.scala 67:65]
    end
    if (reset) begin // @[H2C.scala 29:42]
      send_cmd_count <= 32'h0; // @[H2C.scala 29:42]
    end else if (_T_2) begin // @[H2C.scala 84:32]
      send_cmd_count <= _send_cmd_count_T_1; // @[H2C.scala 85:33]
    end
    complete <= reset | _GEN_21; // @[H2C.scala 32:42 H2C.scala 32:42]
    if (reset) begin // @[H2C.scala 34:50]
      hold <= 4'h0; // @[H2C.scala 34:50]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[H2C.scala 69:48]
          hold <= 4'ha; // @[H2C.scala 72:65]
        end
      end else if (_T_3) begin // @[Conditional.scala 39:67]
        hold <= _hold_T_1; // @[H2C.scala 76:30]
      end
    end
    if (reset) begin // @[H2C.scala 52:42]
      state_cmd <= 2'h0; // @[H2C.scala 52:42]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2C.scala 56:39]
        state_cmd <= 2'h1; // @[H2C.scala 57:65]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (_T_2) begin // @[H2C.scala 69:48]
        state_cmd <= 2'h2; // @[H2C.scala 70:65]
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      state_cmd <= _GEN_11;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  length = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  valid_cmd = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  count_time = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  send_cmd_count = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  complete = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  hold = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  state_cmd = _RAND_7[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue_18(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_c2h_start_addr,
  input  [33:0] io_in_bits_m2h_start_addr,
  input  [31:0] io_in_bits_m2h_length,
  input  [63:0] io_in_bits_c2h_cpt_addr,
  input  [31:0] io_in_bits_pkt_size,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_c2h_start_addr,
  output [33:0] io_out_bits_m2h_start_addr,
  output [31:0] io_out_bits_m2h_length,
  output [63:0] io_out_bits_c2h_cpt_addr,
  output [31:0] io_out_bits_pkt_size
);
  wire  fifo_io_m_clk; // @[XQueue.scala 67:42]
  wire  fifo_io_s_clk; // @[XQueue.scala 67:42]
  wire  fifo_io_reset_n; // @[XQueue.scala 67:42]
  wire [231:0] fifo_io_in_data; // @[XQueue.scala 67:42]
  wire  fifo_io_in_valid; // @[XQueue.scala 67:42]
  wire [231:0] fifo_io_out_data; // @[XQueue.scala 67:42]
  wire  fifo_io_out_valid; // @[XQueue.scala 67:42]
  wire  fifo_io_out_ready; // @[XQueue.scala 67:42]
  wire [225:0] _fifo_io_in_data_T = {io_in_bits_c2h_start_addr,io_in_bits_m2h_start_addr,io_in_bits_m2h_length,
    io_in_bits_c2h_cpt_addr,io_in_bits_pkt_size}; // @[XQueue.scala 73:71]
  SV_STREAM_FIFO_5 fifo ( // @[XQueue.scala 67:42]
    .io_m_clk(fifo_io_m_clk),
    .io_s_clk(fifo_io_s_clk),
    .io_reset_n(fifo_io_reset_n),
    .io_in_data(fifo_io_in_data),
    .io_in_valid(fifo_io_in_valid),
    .io_out_data(fifo_io_out_data),
    .io_out_valid(fifo_io_out_valid),
    .io_out_ready(fifo_io_out_ready)
  );
  assign io_out_valid = fifo_io_out_valid; // @[XQueue.scala 78:49]
  assign io_out_bits_c2h_start_addr = fifo_io_out_data[225:162]; // @[XQueue.scala 77:85]
  assign io_out_bits_m2h_start_addr = fifo_io_out_data[161:128]; // @[XQueue.scala 77:85]
  assign io_out_bits_m2h_length = fifo_io_out_data[127:96]; // @[XQueue.scala 77:85]
  assign io_out_bits_c2h_cpt_addr = fifo_io_out_data[95:32]; // @[XQueue.scala 77:85]
  assign io_out_bits_pkt_size = fifo_io_out_data[31:0]; // @[XQueue.scala 77:85]
  assign fifo_io_m_clk = clock; // @[XQueue.scala 70:49]
  assign fifo_io_s_clk = clock; // @[XQueue.scala 69:49]
  assign fifo_io_reset_n = ~reset; // @[XQueue.scala 71:52]
  assign fifo_io_in_data = {{6'd0}, _fifo_io_in_data_T}; // @[XQueue.scala 73:71]
  assign fifo_io_in_valid = io_in_valid; // @[XQueue.scala 74:49]
  assign fifo_io_out_ready = io_out_ready; // @[XQueue.scala 79:49]
endmodule
module d2hcmdqueuehead(
  input         clock,
  input         reset,
  output        io_cmd_in_ready,
  input         io_cmd_in_valid,
  input  [63:0] io_cmd_in_bits_c2h_start_addr,
  input  [33:0] io_cmd_in_bits_m2h_start_addr,
  input  [31:0] io_cmd_in_bits_m2h_length,
  input  [63:0] io_cmd_in_bits_c2h_cpt_addr,
  input  [31:0] io_cmd_in_bits_pkt_size,
  input         io_cmd_out_ready,
  output        io_cmd_out_valid,
  output [63:0] io_cmd_out_bits_c2h_start_addr,
  output [33:0] io_cmd_out_bits_m2h_start_addr,
  output [31:0] io_cmd_out_bits_m2h_length,
  output [63:0] io_cmd_out_bits_c2h_cpt_addr,
  output [31:0] io_c2h_length,
  output        io_m2h_complete,
  input         io_c2h_finish,
  input         io_m2h_finish,
  input         io_m2h_cpt_complete,
  output        io_last,
  output        io_working,
  output        io_continue
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg  cmd_in_ready; // @[d2hcmdqueuehead.scala 24:46]
  reg  cmd_out_valid; // @[d2hcmdqueuehead.scala 25:46]
  reg  m2h_complete; // @[d2hcmdqueuehead.scala 26:46]
  reg  working; // @[d2hcmdqueuehead.scala 27:46]
  reg  last; // @[d2hcmdqueuehead.scala 28:46]
  reg  continue_; // @[d2hcmdqueuehead.scala 29:46]
  reg [31:0] length; // @[d2hcmdqueuehead.scala 37:46]
  reg [63:0] c2h_addr; // @[d2hcmdqueuehead.scala 38:46]
  reg [33:0] m2h_addr; // @[d2hcmdqueuehead.scala 39:46]
  reg [31:0] length_reg; // @[d2hcmdqueuehead.scala 40:46]
  reg [33:0] m2h_addr_reg; // @[d2hcmdqueuehead.scala 41:46]
  reg [33:0] next_addr; // @[d2hcmdqueuehead.scala 42:46]
  reg [33:0] end_addr; // @[d2hcmdqueuehead.scala 43:46]
  reg [63:0] c2h_cpt_addr; // @[d2hcmdqueuehead.scala 44:46]
  reg [31:0] pkt_size; // @[d2hcmdqueuehead.scala 45:46]
  wire  _T = io_cmd_in_ready & io_cmd_in_valid; // @[Decoupled.scala 40:37]
  wire [33:0] _GEN_39 = {{2'd0}, io_cmd_in_bits_m2h_length}; // @[d2hcmdqueuehead.scala 64:70]
  wire [33:0] _end_addr_T_1 = io_cmd_in_bits_m2h_start_addr + _GEN_39; // @[d2hcmdqueuehead.scala 64:70]
  wire [33:0] _GEN_40 = {{2'd0}, io_cmd_in_bits_pkt_size}; // @[d2hcmdqueuehead.scala 73:70]
  wire [33:0] _next_addr_T_1 = io_cmd_in_bits_m2h_start_addr + _GEN_40; // @[d2hcmdqueuehead.scala 73:70]
  wire [31:0] _GEN_0 = io_cmd_in_bits_m2h_length > io_cmd_in_bits_pkt_size ? io_cmd_in_bits_pkt_size :
    io_cmd_in_bits_m2h_length; // @[d2hcmdqueuehead.scala 70:67 d2hcmdqueuehead.scala 71:37 d2hcmdqueuehead.scala 75:37]
  wire [33:0] _GEN_1 = io_cmd_in_bits_m2h_length > io_cmd_in_bits_pkt_size ? _next_addr_T_1 : _end_addr_T_1; // @[d2hcmdqueuehead.scala 70:67 d2hcmdqueuehead.scala 73:37 d2hcmdqueuehead.scala 77:37]
  wire [63:0] _GEN_2 = _T ? io_cmd_in_bits_c2h_start_addr : c2h_addr; // @[d2hcmdqueuehead.scala 60:27 d2hcmdqueuehead.scala 61:37 d2hcmdqueuehead.scala 38:46]
  wire [33:0] _GEN_3 = _T ? io_cmd_in_bits_m2h_start_addr : m2h_addr; // @[d2hcmdqueuehead.scala 60:27 d2hcmdqueuehead.scala 62:37 d2hcmdqueuehead.scala 39:46]
  wire [31:0] _GEN_8 = _T ? _GEN_0 : length; // @[d2hcmdqueuehead.scala 60:27 d2hcmdqueuehead.scala 37:46]
  wire [33:0] _GEN_10 = _T ? _GEN_1 : next_addr; // @[d2hcmdqueuehead.scala 60:27 d2hcmdqueuehead.scala 42:46]
  wire  _GEN_11 = _T ? 1'h0 : cmd_in_ready; // @[d2hcmdqueuehead.scala 60:27 d2hcmdqueuehead.scala 79:37 d2hcmdqueuehead.scala 24:46]
  wire  _GEN_12 = _T | cmd_out_valid; // @[d2hcmdqueuehead.scala 60:27 d2hcmdqueuehead.scala 80:37 d2hcmdqueuehead.scala 25:46]
  wire  _GEN_13 = _T | working; // @[d2hcmdqueuehead.scala 60:27 d2hcmdqueuehead.scala 81:37 d2hcmdqueuehead.scala 27:46]
  wire  _T_2 = io_cmd_out_ready & io_cmd_out_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_42 = {{32'd0}, length}; // @[d2hcmdqueuehead.scala 93:49]
  wire [63:0] _c2h_addr_T_1 = c2h_addr + _GEN_42; // @[d2hcmdqueuehead.scala 93:49]
  wire [33:0] _GEN_43 = {{2'd0}, length}; // @[d2hcmdqueuehead.scala 94:49]
  wire [33:0] _m2h_addr_T_1 = m2h_addr + _GEN_43; // @[d2hcmdqueuehead.scala 94:49]
  wire [33:0] _T_5 = next_addr + _GEN_43; // @[d2hcmdqueuehead.scala 95:29]
  wire [33:0] _length_T_1 = end_addr - next_addr; // @[d2hcmdqueuehead.scala 99:49]
  wire [33:0] _GEN_14 = _T_5 < end_addr ? {{2'd0}, pkt_size} : _length_T_1; // @[d2hcmdqueuehead.scala 95:49 d2hcmdqueuehead.scala 96:37 d2hcmdqueuehead.scala 99:37]
  wire  _GEN_17 = next_addr == end_addr | last; // @[d2hcmdqueuehead.scala 87:38 d2hcmdqueuehead.scala 89:37 d2hcmdqueuehead.scala 28:46]
  wire  _GEN_18 = next_addr == end_addr ? 1'h0 : 1'h1; // @[d2hcmdqueuehead.scala 87:38 d2hcmdqueuehead.scala 90:37 d2hcmdqueuehead.scala 92:37]
  wire [33:0] _GEN_21 = next_addr == end_addr ? {{2'd0}, _GEN_8} : _GEN_14; // @[d2hcmdqueuehead.scala 87:38]
  wire  _GEN_27 = _T_2 ? _GEN_18 : continue_; // @[d2hcmdqueuehead.scala 84:28 d2hcmdqueuehead.scala 29:46]
  wire [33:0] _GEN_30 = _T_2 ? _GEN_21 : {{2'd0}, _GEN_8}; // @[d2hcmdqueuehead.scala 84:28]
  wire  _GEN_32 = continue_ ? 1'h0 : _GEN_27; // @[d2hcmdqueuehead.scala 105:20 d2hcmdqueuehead.scala 106:25]
  wire  _GEN_33 = last & io_c2h_finish & io_m2h_finish | m2h_complete; // @[d2hcmdqueuehead.scala 109:48 d2hcmdqueuehead.scala 110:25 d2hcmdqueuehead.scala 26:46]
  wire  _GEN_36 = last & m2h_complete & io_m2h_cpt_complete | _GEN_11; // @[d2hcmdqueuehead.scala 113:53 d2hcmdqueuehead.scala 116:25]
  wire  _GEN_38 = last & m2h_complete & io_m2h_cpt_complete | _GEN_32; // @[d2hcmdqueuehead.scala 113:53 d2hcmdqueuehead.scala 118:25]
  assign io_cmd_in_ready = cmd_in_ready; // @[d2hcmdqueuehead.scala 30:37]
  assign io_cmd_out_valid = cmd_out_valid; // @[d2hcmdqueuehead.scala 31:37]
  assign io_cmd_out_bits_c2h_start_addr = c2h_addr; // @[d2hcmdqueuehead.scala 51:37]
  assign io_cmd_out_bits_m2h_start_addr = m2h_addr_reg; // @[d2hcmdqueuehead.scala 52:37]
  assign io_cmd_out_bits_m2h_length = length_reg; // @[d2hcmdqueuehead.scala 49:37]
  assign io_cmd_out_bits_c2h_cpt_addr = c2h_cpt_addr; // @[d2hcmdqueuehead.scala 57:37]
  assign io_c2h_length = length; // @[d2hcmdqueuehead.scala 50:37]
  assign io_m2h_complete = m2h_complete; // @[d2hcmdqueuehead.scala 32:37]
  assign io_last = last; // @[d2hcmdqueuehead.scala 33:37]
  assign io_working = working; // @[d2hcmdqueuehead.scala 34:37]
  assign io_continue = continue_; // @[d2hcmdqueuehead.scala 35:37]
  always @(posedge clock) begin
    cmd_in_ready <= reset | _GEN_36; // @[d2hcmdqueuehead.scala 24:46 d2hcmdqueuehead.scala 24:46]
    if (reset) begin // @[d2hcmdqueuehead.scala 25:46]
      cmd_out_valid <= 1'h0; // @[d2hcmdqueuehead.scala 25:46]
    end else if (_T_2) begin // @[d2hcmdqueuehead.scala 84:28]
      if (next_addr == end_addr) begin // @[d2hcmdqueuehead.scala 87:38]
        cmd_out_valid <= 1'h0; // @[d2hcmdqueuehead.scala 88:37]
      end else begin
        cmd_out_valid <= _GEN_12;
      end
    end else begin
      cmd_out_valid <= _GEN_12;
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 26:46]
      m2h_complete <= 1'h0; // @[d2hcmdqueuehead.scala 26:46]
    end else if (last & m2h_complete & io_m2h_cpt_complete) begin // @[d2hcmdqueuehead.scala 113:53]
      m2h_complete <= 1'h0; // @[d2hcmdqueuehead.scala 114:25]
    end else begin
      m2h_complete <= _GEN_33;
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 27:46]
      working <= 1'h0; // @[d2hcmdqueuehead.scala 27:46]
    end else if (last & m2h_complete & io_m2h_cpt_complete) begin // @[d2hcmdqueuehead.scala 113:53]
      working <= 1'h0; // @[d2hcmdqueuehead.scala 117:25]
    end else begin
      working <= _GEN_13;
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 28:46]
      last <= 1'h0; // @[d2hcmdqueuehead.scala 28:46]
    end else if (last & m2h_complete & io_m2h_cpt_complete) begin // @[d2hcmdqueuehead.scala 113:53]
      last <= 1'h0; // @[d2hcmdqueuehead.scala 115:25]
    end else if (_T_2) begin // @[d2hcmdqueuehead.scala 84:28]
      last <= _GEN_17;
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 29:46]
      continue_ <= 1'h0; // @[d2hcmdqueuehead.scala 29:46]
    end else begin
      continue_ <= _GEN_38;
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 37:46]
      length <= 32'h0; // @[d2hcmdqueuehead.scala 37:46]
    end else begin
      length <= _GEN_30[31:0];
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 38:46]
      c2h_addr <= 64'h0; // @[d2hcmdqueuehead.scala 38:46]
    end else if (_T_2) begin // @[d2hcmdqueuehead.scala 84:28]
      if (next_addr == end_addr) begin // @[d2hcmdqueuehead.scala 87:38]
        c2h_addr <= _GEN_2;
      end else begin
        c2h_addr <= _c2h_addr_T_1; // @[d2hcmdqueuehead.scala 93:37]
      end
    end else begin
      c2h_addr <= _GEN_2;
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 39:46]
      m2h_addr <= 34'h0; // @[d2hcmdqueuehead.scala 39:46]
    end else if (_T_2) begin // @[d2hcmdqueuehead.scala 84:28]
      if (next_addr == end_addr) begin // @[d2hcmdqueuehead.scala 87:38]
        m2h_addr <= _GEN_3;
      end else begin
        m2h_addr <= _m2h_addr_T_1; // @[d2hcmdqueuehead.scala 94:37]
      end
    end else begin
      m2h_addr <= _GEN_3;
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 40:46]
      length_reg <= 32'h0; // @[d2hcmdqueuehead.scala 40:46]
    end else if (_T_2) begin // @[d2hcmdqueuehead.scala 84:28]
      length_reg <= length; // @[d2hcmdqueuehead.scala 85:37]
    end else if (_T) begin // @[d2hcmdqueuehead.scala 60:27]
      if (io_cmd_in_bits_m2h_length > io_cmd_in_bits_pkt_size) begin // @[d2hcmdqueuehead.scala 70:67]
        length_reg <= io_cmd_in_bits_pkt_size; // @[d2hcmdqueuehead.scala 71:37]
      end else begin
        length_reg <= io_cmd_in_bits_m2h_length; // @[d2hcmdqueuehead.scala 75:37]
      end
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 41:46]
      m2h_addr_reg <= 34'h0; // @[d2hcmdqueuehead.scala 41:46]
    end else if (_T_2) begin // @[d2hcmdqueuehead.scala 84:28]
      m2h_addr_reg <= m2h_addr; // @[d2hcmdqueuehead.scala 86:37]
    end else if (_T) begin // @[d2hcmdqueuehead.scala 60:27]
      m2h_addr_reg <= io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueuehead.scala 63:37]
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 42:46]
      next_addr <= 34'h0; // @[d2hcmdqueuehead.scala 42:46]
    end else if (_T_2) begin // @[d2hcmdqueuehead.scala 84:28]
      if (next_addr == end_addr) begin // @[d2hcmdqueuehead.scala 87:38]
        next_addr <= _GEN_10;
      end else if (_T_5 < end_addr) begin // @[d2hcmdqueuehead.scala 95:49]
        next_addr <= _T_5; // @[d2hcmdqueuehead.scala 97:37]
      end else begin
        next_addr <= end_addr; // @[d2hcmdqueuehead.scala 100:37]
      end
    end else begin
      next_addr <= _GEN_10;
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 43:46]
      end_addr <= 34'h0; // @[d2hcmdqueuehead.scala 43:46]
    end else if (_T) begin // @[d2hcmdqueuehead.scala 60:27]
      end_addr <= _end_addr_T_1; // @[d2hcmdqueuehead.scala 64:37]
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 44:46]
      c2h_cpt_addr <= 64'h0; // @[d2hcmdqueuehead.scala 44:46]
    end else if (_T) begin // @[d2hcmdqueuehead.scala 60:27]
      c2h_cpt_addr <= io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueuehead.scala 65:37]
    end
    if (reset) begin // @[d2hcmdqueuehead.scala 45:46]
      pkt_size <= 32'h1000; // @[d2hcmdqueuehead.scala 45:46]
    end else if (_T) begin // @[d2hcmdqueuehead.scala 60:27]
      pkt_size <= io_cmd_in_bits_pkt_size; // @[d2hcmdqueuehead.scala 66:37]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cmd_in_ready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cmd_out_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  m2h_complete = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  working = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  last = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  continue_ = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  length = _RAND_6[31:0];
  _RAND_7 = {2{`RANDOM}};
  c2h_addr = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  m2h_addr = _RAND_8[33:0];
  _RAND_9 = {1{`RANDOM}};
  length_reg = _RAND_9[31:0];
  _RAND_10 = {2{`RANDOM}};
  m2h_addr_reg = _RAND_10[33:0];
  _RAND_11 = {2{`RANDOM}};
  next_addr = _RAND_11[33:0];
  _RAND_12 = {2{`RANDOM}};
  end_addr = _RAND_12[33:0];
  _RAND_13 = {2{`RANDOM}};
  c2h_cpt_addr = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  pkt_size = _RAND_14[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module d2hcmdqueue(
  input         clock,
  input         reset,
  input         io_cmd_in_valid,
  input  [63:0] io_cmd_in_bits_c2h_start_addr,
  input  [33:0] io_cmd_in_bits_m2h_start_addr,
  input  [31:0] io_cmd_in_bits_m2h_length,
  input  [63:0] io_cmd_in_bits_c2h_cpt_addr,
  input  [31:0] io_cmd_in_bits_pkt_size,
  input  [31:0] io_qin,
  input         io_cmd_out_ready,
  output        io_cmd_out_valid,
  output [63:0] io_cmd_out_bits_c2h_start_addr,
  output [33:0] io_cmd_out_bits_m2h_start_addr,
  output [31:0] io_cmd_out_bits_m2h_length,
  output [63:0] io_cmd_out_bits_c2h_cpt_addr,
  output [31:0] io_c2h_length,
  output        io_m2h_complete,
  input         io_c2h_finish,
  input         io_m2h_finish,
  input         io_m2h_cpt_complete,
  input         io_read_count_equal,
  input         io_empty,
  input         io_h2m_complete_start,
  output        io_h2m_complete,
  input         io_h2m_cpt_complete,
  input         io_m2h_valid_tmpreg,
  output        io_last,
  output [31:0] io_counter
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  Q_0_clock; // @[XQueue.scala 35:23]
  wire  Q_0_reset; // @[XQueue.scala 35:23]
  wire  Q_0_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_0_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_0_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_0_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_0_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_0_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_0_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_0_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_0_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_0_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_0_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_0_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_0_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_1_clock; // @[XQueue.scala 35:23]
  wire  Q_1_reset; // @[XQueue.scala 35:23]
  wire  Q_1_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_1_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_1_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_1_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_1_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_1_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_1_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_1_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_1_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_1_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_1_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_1_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_1_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_2_clock; // @[XQueue.scala 35:23]
  wire  Q_2_reset; // @[XQueue.scala 35:23]
  wire  Q_2_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_2_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_2_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_2_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_2_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_2_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_2_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_2_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_2_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_2_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_2_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_2_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_2_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_3_clock; // @[XQueue.scala 35:23]
  wire  Q_3_reset; // @[XQueue.scala 35:23]
  wire  Q_3_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_3_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_3_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_3_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_3_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_3_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_3_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_3_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_3_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_3_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_3_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_3_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_3_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_4_clock; // @[XQueue.scala 35:23]
  wire  Q_4_reset; // @[XQueue.scala 35:23]
  wire  Q_4_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_4_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_4_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_4_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_4_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_4_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_4_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_4_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_4_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_4_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_4_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_4_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_4_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_5_clock; // @[XQueue.scala 35:23]
  wire  Q_5_reset; // @[XQueue.scala 35:23]
  wire  Q_5_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_5_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_5_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_5_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_5_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_5_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_5_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_5_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_5_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_5_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_5_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_5_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_5_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_6_clock; // @[XQueue.scala 35:23]
  wire  Q_6_reset; // @[XQueue.scala 35:23]
  wire  Q_6_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_6_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_6_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_6_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_6_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_6_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_6_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_6_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_6_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_6_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_6_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_6_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_6_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_7_clock; // @[XQueue.scala 35:23]
  wire  Q_7_reset; // @[XQueue.scala 35:23]
  wire  Q_7_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_7_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_7_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_7_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_7_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_7_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_7_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_7_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_7_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_7_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_7_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_7_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_7_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_8_clock; // @[XQueue.scala 35:23]
  wire  Q_8_reset; // @[XQueue.scala 35:23]
  wire  Q_8_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_8_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_8_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_8_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_8_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_8_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_8_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_8_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_8_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_8_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_8_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_8_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_8_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_9_clock; // @[XQueue.scala 35:23]
  wire  Q_9_reset; // @[XQueue.scala 35:23]
  wire  Q_9_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_9_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_9_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_9_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_9_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_9_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_9_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_9_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_9_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_9_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_9_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_9_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_9_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_10_clock; // @[XQueue.scala 35:23]
  wire  Q_10_reset; // @[XQueue.scala 35:23]
  wire  Q_10_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_10_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_10_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_10_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_10_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_10_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_10_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_10_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_10_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_10_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_10_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_10_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_10_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_11_clock; // @[XQueue.scala 35:23]
  wire  Q_11_reset; // @[XQueue.scala 35:23]
  wire  Q_11_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_11_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_11_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_11_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_11_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_11_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_11_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_11_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_11_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_11_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_11_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_11_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_11_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_12_clock; // @[XQueue.scala 35:23]
  wire  Q_12_reset; // @[XQueue.scala 35:23]
  wire  Q_12_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_12_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_12_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_12_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_12_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_12_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_12_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_12_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_12_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_12_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_12_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_12_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_12_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_13_clock; // @[XQueue.scala 35:23]
  wire  Q_13_reset; // @[XQueue.scala 35:23]
  wire  Q_13_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_13_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_13_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_13_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_13_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_13_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_13_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_13_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_13_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_13_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_13_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_13_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_13_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_14_clock; // @[XQueue.scala 35:23]
  wire  Q_14_reset; // @[XQueue.scala 35:23]
  wire  Q_14_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_14_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_14_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_14_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_14_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_14_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_14_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_14_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_14_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_14_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_14_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_14_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_14_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_15_clock; // @[XQueue.scala 35:23]
  wire  Q_15_reset; // @[XQueue.scala 35:23]
  wire  Q_15_io_in_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_15_io_in_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_15_io_in_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_15_io_in_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_15_io_in_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_15_io_in_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Q_15_io_out_ready; // @[XQueue.scala 35:23]
  wire  Q_15_io_out_valid; // @[XQueue.scala 35:23]
  wire [63:0] Q_15_io_out_bits_c2h_start_addr; // @[XQueue.scala 35:23]
  wire [33:0] Q_15_io_out_bits_m2h_start_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_15_io_out_bits_m2h_length; // @[XQueue.scala 35:23]
  wire [63:0] Q_15_io_out_bits_c2h_cpt_addr; // @[XQueue.scala 35:23]
  wire [31:0] Q_15_io_out_bits_pkt_size; // @[XQueue.scala 35:23]
  wire  Qh_0_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_0_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_0_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_0_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_0_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_0_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_0_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_0_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_0_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_0_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_0_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_0_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_1_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_1_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_1_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_1_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_1_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_1_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_1_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_1_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_1_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_1_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_1_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_2_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_2_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_2_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_2_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_2_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_2_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_2_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_2_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_2_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_2_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_2_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_3_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_3_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_3_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_3_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_3_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_3_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_3_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_3_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_3_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_3_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_3_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_4_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_4_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_4_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_4_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_4_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_4_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_4_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_4_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_4_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_4_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_4_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_5_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_5_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_5_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_5_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_5_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_5_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_5_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_5_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_5_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_5_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_5_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_6_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_6_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_6_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_6_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_6_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_6_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_6_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_6_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_6_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_6_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_6_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_7_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_7_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_7_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_7_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_7_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_7_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_7_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_7_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_7_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_7_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_7_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_8_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_8_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_8_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_8_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_8_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_8_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_8_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_8_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_8_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_8_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_8_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_9_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_9_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_9_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_9_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_9_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_9_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_9_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_9_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_9_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_9_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_9_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_10_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_10_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_10_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_10_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_10_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_10_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_10_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_10_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_10_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_10_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_10_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_11_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_11_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_11_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_11_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_11_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_11_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_11_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_11_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_11_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_11_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_11_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_12_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_12_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_12_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_12_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_12_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_12_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_12_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_12_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_12_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_12_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_12_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_13_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_13_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_13_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_13_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_13_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_13_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_13_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_13_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_13_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_13_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_13_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_14_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_14_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_14_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_14_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_14_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_14_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_14_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_14_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_14_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_14_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_14_io_continue; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_clock; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_reset; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_cmd_in_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_cmd_in_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_15_io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_15_io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_15_io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_15_io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_15_io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_cmd_out_ready; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_cmd_out_valid; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_15_io_cmd_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [33:0] Qh_15_io_cmd_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_15_io_cmd_out_bits_m2h_length; // @[d2hcmdqueue.scala 35:45]
  wire [63:0] Qh_15_io_cmd_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 35:45]
  wire [31:0] Qh_15_io_c2h_length; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_m2h_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_c2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_m2h_finish; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_m2h_cpt_complete; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_last; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_working; // @[d2hcmdqueue.scala 35:45]
  wire  Qh_15_io_continue; // @[d2hcmdqueue.scala 35:45]
  reg [31:0] counter; // @[d2hcmdqueue.scala 37:26]
  wire  _T = io_cmd_out_ready & io_cmd_out_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[d2hcmdqueue.scala 41:28]
  reg  h2m_cpt_working; // @[d2hcmdqueue.scala 46:34]
  reg  h2m_complete; // @[d2hcmdqueue.scala 47:31]
  wire  _GEN_1 = io_h2m_complete_start | h2m_cpt_working; // @[d2hcmdqueue.scala 50:5 d2hcmdqueue.scala 51:25 d2hcmdqueue.scala 46:34]
  reg [4:0] out; // @[d2hcmdqueue.scala 54:23]
  reg [4:0] next; // @[d2hcmdqueue.scala 55:23]
  reg [4:0] hold1; // @[d2hcmdqueue.scala 56:24]
  reg [4:0] hold2; // @[d2hcmdqueue.scala 57:24]
  wire  _Qh_0_io_cmd_out_ready_T = out == 5'h0; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_1_io_cmd_out_ready_T = out == 5'h1; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_2_io_cmd_out_ready_T = out == 5'h2; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_3_io_cmd_out_ready_T = out == 5'h3; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_4_io_cmd_out_ready_T = out == 5'h4; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_5_io_cmd_out_ready_T = out == 5'h5; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_6_io_cmd_out_ready_T = out == 5'h6; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_7_io_cmd_out_ready_T = out == 5'h7; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_8_io_cmd_out_ready_T = out == 5'h8; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_9_io_cmd_out_ready_T = out == 5'h9; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_10_io_cmd_out_ready_T = out == 5'ha; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_11_io_cmd_out_ready_T = out == 5'hb; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_12_io_cmd_out_ready_T = out == 5'hc; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_13_io_cmd_out_ready_T = out == 5'hd; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_14_io_cmd_out_ready_T = out == 5'he; // @[d2hcmdqueue.scala 63:64]
  wire  _Qh_15_io_cmd_out_ready_T = out == 5'hf; // @[d2hcmdqueue.scala 63:64]
  wire  _T_1 = ~Qh_0_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_3 = ~Qh_0_io_working & _Qh_0_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire  _T_4 = ~h2m_cpt_working; // @[d2hcmdqueue.scala 72:60]
  wire [4:0] _GEN_2 = _T_3 & h2m_cpt_working ? 5'h1f : out; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17 d2hcmdqueue.scala 54:23]
  wire [4:0] _GEN_3 = ~Qh_0_io_working & _Qh_0_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_2; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_12 = Qh_0_io_continue & _Qh_0_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _T_16 = 5'h10 - 5'h1; // @[d2hcmdqueue.scala 80:36]
  wire [4:0] _next_T_1 = next + 5'h1; // @[d2hcmdqueue.scala 83:30]
  wire [4:0] _GEN_4 = next == _T_16 ? 5'h0 : _next_T_1; // @[d2hcmdqueue.scala 80:42 d2hcmdqueue.scala 81:22 d2hcmdqueue.scala 83:22]
  wire [4:0] _GEN_5 = _T_12 & h2m_cpt_working ? 5'h1f : _GEN_3; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_6 = Qh_0_io_continue & _Qh_0_io_cmd_out_ready_T & _T_4 ? next : _GEN_5; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_7 = Qh_0_io_continue & _Qh_0_io_cmd_out_ready_T & _T_4 ? _GEN_4 : next; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 55:23]
  wire [4:0] _GEN_9 = _T_1 & next == 5'h0 ? _GEN_4 : _GEN_7; // @[d2hcmdqueue.scala 89:58]
  wire  _T_28 = ~Qh_1_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_30 = ~Qh_1_io_working & _Qh_1_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_10 = _T_30 & h2m_cpt_working ? 5'h1f : _GEN_6; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_11 = ~Qh_1_io_working & _Qh_1_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_10; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_39 = Qh_1_io_continue & _Qh_1_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_13 = _T_39 & h2m_cpt_working ? 5'h1f : _GEN_11; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_14 = Qh_1_io_continue & _Qh_1_io_cmd_out_ready_T & _T_4 ? next : _GEN_13; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_15 = Qh_1_io_continue & _Qh_1_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_9; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_17 = _T_28 & next == 5'h1 ? _GEN_4 : _GEN_15; // @[d2hcmdqueue.scala 89:58]
  wire  _T_55 = ~Qh_2_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_57 = ~Qh_2_io_working & _Qh_2_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_18 = _T_57 & h2m_cpt_working ? 5'h1f : _GEN_14; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_19 = ~Qh_2_io_working & _Qh_2_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_18; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_66 = Qh_2_io_continue & _Qh_2_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_21 = _T_66 & h2m_cpt_working ? 5'h1f : _GEN_19; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_22 = Qh_2_io_continue & _Qh_2_io_cmd_out_ready_T & _T_4 ? next : _GEN_21; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_23 = Qh_2_io_continue & _Qh_2_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_17; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_25 = _T_55 & next == 5'h2 ? _GEN_4 : _GEN_23; // @[d2hcmdqueue.scala 89:58]
  wire  _T_82 = ~Qh_3_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_84 = ~Qh_3_io_working & _Qh_3_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_26 = _T_84 & h2m_cpt_working ? 5'h1f : _GEN_22; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_27 = ~Qh_3_io_working & _Qh_3_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_26; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_93 = Qh_3_io_continue & _Qh_3_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_29 = _T_93 & h2m_cpt_working ? 5'h1f : _GEN_27; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_30 = Qh_3_io_continue & _Qh_3_io_cmd_out_ready_T & _T_4 ? next : _GEN_29; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_31 = Qh_3_io_continue & _Qh_3_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_25; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_33 = _T_82 & next == 5'h3 ? _GEN_4 : _GEN_31; // @[d2hcmdqueue.scala 89:58]
  wire  _T_109 = ~Qh_4_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_111 = ~Qh_4_io_working & _Qh_4_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_34 = _T_111 & h2m_cpt_working ? 5'h1f : _GEN_30; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_35 = ~Qh_4_io_working & _Qh_4_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_34; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_120 = Qh_4_io_continue & _Qh_4_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_37 = _T_120 & h2m_cpt_working ? 5'h1f : _GEN_35; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_38 = Qh_4_io_continue & _Qh_4_io_cmd_out_ready_T & _T_4 ? next : _GEN_37; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_39 = Qh_4_io_continue & _Qh_4_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_33; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_41 = _T_109 & next == 5'h4 ? _GEN_4 : _GEN_39; // @[d2hcmdqueue.scala 89:58]
  wire  _T_136 = ~Qh_5_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_138 = ~Qh_5_io_working & _Qh_5_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_42 = _T_138 & h2m_cpt_working ? 5'h1f : _GEN_38; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_43 = ~Qh_5_io_working & _Qh_5_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_42; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_147 = Qh_5_io_continue & _Qh_5_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_45 = _T_147 & h2m_cpt_working ? 5'h1f : _GEN_43; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_46 = Qh_5_io_continue & _Qh_5_io_cmd_out_ready_T & _T_4 ? next : _GEN_45; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_47 = Qh_5_io_continue & _Qh_5_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_41; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_49 = _T_136 & next == 5'h5 ? _GEN_4 : _GEN_47; // @[d2hcmdqueue.scala 89:58]
  wire  _T_163 = ~Qh_6_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_165 = ~Qh_6_io_working & _Qh_6_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_50 = _T_165 & h2m_cpt_working ? 5'h1f : _GEN_46; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_51 = ~Qh_6_io_working & _Qh_6_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_50; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_174 = Qh_6_io_continue & _Qh_6_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_53 = _T_174 & h2m_cpt_working ? 5'h1f : _GEN_51; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_54 = Qh_6_io_continue & _Qh_6_io_cmd_out_ready_T & _T_4 ? next : _GEN_53; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_55 = Qh_6_io_continue & _Qh_6_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_49; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_57 = _T_163 & next == 5'h6 ? _GEN_4 : _GEN_55; // @[d2hcmdqueue.scala 89:58]
  wire  _T_190 = ~Qh_7_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_192 = ~Qh_7_io_working & _Qh_7_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_58 = _T_192 & h2m_cpt_working ? 5'h1f : _GEN_54; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_59 = ~Qh_7_io_working & _Qh_7_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_58; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_201 = Qh_7_io_continue & _Qh_7_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_61 = _T_201 & h2m_cpt_working ? 5'h1f : _GEN_59; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_62 = Qh_7_io_continue & _Qh_7_io_cmd_out_ready_T & _T_4 ? next : _GEN_61; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_63 = Qh_7_io_continue & _Qh_7_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_57; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_65 = _T_190 & next == 5'h7 ? _GEN_4 : _GEN_63; // @[d2hcmdqueue.scala 89:58]
  wire  _T_217 = ~Qh_8_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_219 = ~Qh_8_io_working & _Qh_8_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_66 = _T_219 & h2m_cpt_working ? 5'h1f : _GEN_62; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_67 = ~Qh_8_io_working & _Qh_8_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_66; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_228 = Qh_8_io_continue & _Qh_8_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_69 = _T_228 & h2m_cpt_working ? 5'h1f : _GEN_67; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_70 = Qh_8_io_continue & _Qh_8_io_cmd_out_ready_T & _T_4 ? next : _GEN_69; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_71 = Qh_8_io_continue & _Qh_8_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_65; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_73 = _T_217 & next == 5'h8 ? _GEN_4 : _GEN_71; // @[d2hcmdqueue.scala 89:58]
  wire  _T_244 = ~Qh_9_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_246 = ~Qh_9_io_working & _Qh_9_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_74 = _T_246 & h2m_cpt_working ? 5'h1f : _GEN_70; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_75 = ~Qh_9_io_working & _Qh_9_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_74; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_255 = Qh_9_io_continue & _Qh_9_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_77 = _T_255 & h2m_cpt_working ? 5'h1f : _GEN_75; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_78 = Qh_9_io_continue & _Qh_9_io_cmd_out_ready_T & _T_4 ? next : _GEN_77; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_79 = Qh_9_io_continue & _Qh_9_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_73; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_81 = _T_244 & next == 5'h9 ? _GEN_4 : _GEN_79; // @[d2hcmdqueue.scala 89:58]
  wire  _T_271 = ~Qh_10_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_273 = ~Qh_10_io_working & _Qh_10_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_82 = _T_273 & h2m_cpt_working ? 5'h1f : _GEN_78; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_83 = ~Qh_10_io_working & _Qh_10_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_82; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_282 = Qh_10_io_continue & _Qh_10_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_85 = _T_282 & h2m_cpt_working ? 5'h1f : _GEN_83; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_86 = Qh_10_io_continue & _Qh_10_io_cmd_out_ready_T & _T_4 ? next : _GEN_85; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_87 = Qh_10_io_continue & _Qh_10_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_81; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_89 = _T_271 & next == 5'ha ? _GEN_4 : _GEN_87; // @[d2hcmdqueue.scala 89:58]
  wire  _T_298 = ~Qh_11_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_300 = ~Qh_11_io_working & _Qh_11_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_90 = _T_300 & h2m_cpt_working ? 5'h1f : _GEN_86; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_91 = ~Qh_11_io_working & _Qh_11_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_90; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_309 = Qh_11_io_continue & _Qh_11_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_93 = _T_309 & h2m_cpt_working ? 5'h1f : _GEN_91; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_94 = Qh_11_io_continue & _Qh_11_io_cmd_out_ready_T & _T_4 ? next : _GEN_93; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_95 = Qh_11_io_continue & _Qh_11_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_89; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_97 = _T_298 & next == 5'hb ? _GEN_4 : _GEN_95; // @[d2hcmdqueue.scala 89:58]
  wire  _T_325 = ~Qh_12_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_327 = ~Qh_12_io_working & _Qh_12_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_98 = _T_327 & h2m_cpt_working ? 5'h1f : _GEN_94; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_99 = ~Qh_12_io_working & _Qh_12_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_98; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_336 = Qh_12_io_continue & _Qh_12_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_101 = _T_336 & h2m_cpt_working ? 5'h1f : _GEN_99; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_102 = Qh_12_io_continue & _Qh_12_io_cmd_out_ready_T & _T_4 ? next : _GEN_101; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_103 = Qh_12_io_continue & _Qh_12_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_97; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_105 = _T_325 & next == 5'hc ? _GEN_4 : _GEN_103; // @[d2hcmdqueue.scala 89:58]
  wire  _T_352 = ~Qh_13_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_354 = ~Qh_13_io_working & _Qh_13_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_106 = _T_354 & h2m_cpt_working ? 5'h1f : _GEN_102; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_107 = ~Qh_13_io_working & _Qh_13_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_106; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_363 = Qh_13_io_continue & _Qh_13_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_109 = _T_363 & h2m_cpt_working ? 5'h1f : _GEN_107; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_110 = Qh_13_io_continue & _Qh_13_io_cmd_out_ready_T & _T_4 ? next : _GEN_109; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_111 = Qh_13_io_continue & _Qh_13_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_105; // @[d2hcmdqueue.scala 78:77]
  wire [4:0] _GEN_113 = _T_352 & next == 5'hd ? _GEN_4 : _GEN_111; // @[d2hcmdqueue.scala 89:58]
  wire  _T_379 = ~Qh_14_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_381 = ~Qh_14_io_working & _Qh_14_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_114 = _T_381 & h2m_cpt_working ? 5'h1f : _GEN_110; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_115 = ~Qh_14_io_working & _Qh_14_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_114; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_390 = Qh_14_io_continue & _Qh_14_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_117 = _T_390 & h2m_cpt_working ? 5'h1f : _GEN_115; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_118 = Qh_14_io_continue & _Qh_14_io_cmd_out_ready_T & _T_4 ? next : _GEN_117; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire [4:0] _GEN_119 = Qh_14_io_continue & _Qh_14_io_cmd_out_ready_T & _T_4 ? _GEN_4 : _GEN_113; // @[d2hcmdqueue.scala 78:77]
  wire  _T_406 = ~Qh_15_io_working; // @[d2hcmdqueue.scala 72:32]
  wire  _T_408 = ~Qh_15_io_working & _Qh_15_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 72:44]
  wire [4:0] _GEN_122 = _T_408 & h2m_cpt_working ? 5'h1f : _GEN_118; // @[d2hcmdqueue.scala 75:80 d2hcmdqueue.scala 76:17]
  wire [4:0] _GEN_123 = ~Qh_15_io_working & _Qh_15_io_cmd_out_ready_T & ~h2m_cpt_working ? next : _GEN_122; // @[d2hcmdqueue.scala 72:77 d2hcmdqueue.scala 73:17]
  wire  _T_417 = Qh_15_io_continue & _Qh_15_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 78:44]
  wire [4:0] _GEN_125 = _T_417 & h2m_cpt_working ? 5'h1f : _GEN_123; // @[d2hcmdqueue.scala 86:80 d2hcmdqueue.scala 87:17]
  wire [4:0] _GEN_126 = Qh_15_io_continue & _Qh_15_io_cmd_out_ready_T & _T_4 ? next : _GEN_125; // @[d2hcmdqueue.scala 78:77 d2hcmdqueue.scala 79:17]
  wire  _T_434 = hold1 != 5'h0; // @[d2hcmdqueue.scala 98:21]
  wire [4:0] _hold1_T_1 = hold1 - 5'h1; // @[d2hcmdqueue.scala 99:29]
  wire  _T_437 = io_c2h_finish & io_m2h_finish & io_read_count_equal & io_empty; // @[d2hcmdqueue.scala 100:71]
  wire [4:0] _hold2_T_1 = hold2 - 5'h1; // @[d2hcmdqueue.scala 102:32]
  wire  _T_440 = hold2 == 5'h0 & ~io_m2h_valid_tmpreg; // @[d2hcmdqueue.scala 103:37]
  wire  _GEN_130 = _T_440 | h2m_complete; // @[d2hcmdqueue.scala 104:21 d2hcmdqueue.scala 104:35 d2hcmdqueue.scala 47:31]
  wire [4:0] _GEN_131 = _T_437 ? _hold2_T_1 : hold2; // @[d2hcmdqueue.scala 101:13 d2hcmdqueue.scala 102:23 d2hcmdqueue.scala 57:24]
  wire  _GEN_132 = _T_437 ? _GEN_130 : h2m_complete; // @[d2hcmdqueue.scala 101:13 d2hcmdqueue.scala 47:31]
  wire  _T_441 = h2m_complete & io_h2m_cpt_complete; // @[d2hcmdqueue.scala 106:28]
  wire [63:0] _io_cmd_out_bits_T_1_c2h_start_addr = Qh_0_io_cmd_out_bits_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_1_m2h_start_addr = Qh_0_io_cmd_out_bits_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_1_m2h_length = Qh_0_io_cmd_out_bits_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_1_c2h_cpt_addr = Qh_0_io_cmd_out_bits_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_3_c2h_start_addr = 5'h1 == out ? Qh_1_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_1_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_3_m2h_start_addr = 5'h1 == out ? Qh_1_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_1_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_3_m2h_length = 5'h1 == out ? Qh_1_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_1_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_3_c2h_cpt_addr = 5'h1 == out ? Qh_1_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_1_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_5_c2h_start_addr = 5'h2 == out ? Qh_2_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_3_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_5_m2h_start_addr = 5'h2 == out ? Qh_2_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_3_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_5_m2h_length = 5'h2 == out ? Qh_2_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_3_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_5_c2h_cpt_addr = 5'h2 == out ? Qh_2_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_3_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_7_c2h_start_addr = 5'h3 == out ? Qh_3_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_5_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_7_m2h_start_addr = 5'h3 == out ? Qh_3_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_5_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_7_m2h_length = 5'h3 == out ? Qh_3_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_5_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_7_c2h_cpt_addr = 5'h3 == out ? Qh_3_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_5_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_9_c2h_start_addr = 5'h4 == out ? Qh_4_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_7_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_9_m2h_start_addr = 5'h4 == out ? Qh_4_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_7_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_9_m2h_length = 5'h4 == out ? Qh_4_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_7_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_9_c2h_cpt_addr = 5'h4 == out ? Qh_4_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_7_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_11_c2h_start_addr = 5'h5 == out ? Qh_5_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_9_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_11_m2h_start_addr = 5'h5 == out ? Qh_5_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_9_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_11_m2h_length = 5'h5 == out ? Qh_5_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_9_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_11_c2h_cpt_addr = 5'h5 == out ? Qh_5_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_9_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_13_c2h_start_addr = 5'h6 == out ? Qh_6_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_11_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_13_m2h_start_addr = 5'h6 == out ? Qh_6_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_11_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_13_m2h_length = 5'h6 == out ? Qh_6_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_11_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_13_c2h_cpt_addr = 5'h6 == out ? Qh_6_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_11_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_15_c2h_start_addr = 5'h7 == out ? Qh_7_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_13_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_15_m2h_start_addr = 5'h7 == out ? Qh_7_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_13_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_15_m2h_length = 5'h7 == out ? Qh_7_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_13_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_15_c2h_cpt_addr = 5'h7 == out ? Qh_7_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_13_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_17_c2h_start_addr = 5'h8 == out ? Qh_8_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_15_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_17_m2h_start_addr = 5'h8 == out ? Qh_8_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_15_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_17_m2h_length = 5'h8 == out ? Qh_8_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_15_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_17_c2h_cpt_addr = 5'h8 == out ? Qh_8_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_15_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_19_c2h_start_addr = 5'h9 == out ? Qh_9_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_17_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_19_m2h_start_addr = 5'h9 == out ? Qh_9_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_17_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_19_m2h_length = 5'h9 == out ? Qh_9_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_17_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_19_c2h_cpt_addr = 5'h9 == out ? Qh_9_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_17_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_21_c2h_start_addr = 5'ha == out ? Qh_10_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_19_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_21_m2h_start_addr = 5'ha == out ? Qh_10_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_19_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_21_m2h_length = 5'ha == out ? Qh_10_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_19_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_21_c2h_cpt_addr = 5'ha == out ? Qh_10_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_19_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_23_c2h_start_addr = 5'hb == out ? Qh_11_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_21_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_23_m2h_start_addr = 5'hb == out ? Qh_11_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_21_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_23_m2h_length = 5'hb == out ? Qh_11_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_21_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_23_c2h_cpt_addr = 5'hb == out ? Qh_11_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_21_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_25_c2h_start_addr = 5'hc == out ? Qh_12_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_23_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_25_m2h_start_addr = 5'hc == out ? Qh_12_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_23_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_25_m2h_length = 5'hc == out ? Qh_12_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_23_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_25_c2h_cpt_addr = 5'hc == out ? Qh_12_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_23_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_27_c2h_start_addr = 5'hd == out ? Qh_13_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_25_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_27_m2h_start_addr = 5'hd == out ? Qh_13_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_25_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_27_m2h_length = 5'hd == out ? Qh_13_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_25_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_27_c2h_cpt_addr = 5'hd == out ? Qh_13_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_25_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_29_c2h_start_addr = 5'he == out ? Qh_14_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_27_c2h_start_addr; // @[Mux.scala 80:57]
  wire [33:0] _io_cmd_out_bits_T_29_m2h_start_addr = 5'he == out ? Qh_14_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_27_m2h_start_addr; // @[Mux.scala 80:57]
  wire [31:0] _io_cmd_out_bits_T_29_m2h_length = 5'he == out ? Qh_14_io_cmd_out_bits_m2h_length :
    _io_cmd_out_bits_T_27_m2h_length; // @[Mux.scala 80:57]
  wire [63:0] _io_cmd_out_bits_T_29_c2h_cpt_addr = 5'he == out ? Qh_14_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_27_c2h_cpt_addr; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_3 = 5'h1 == out ? Qh_1_io_cmd_out_valid : Qh_0_io_cmd_out_valid; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_5 = 5'h2 == out ? Qh_2_io_cmd_out_valid : _io_cmd_out_valid_T_3; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_7 = 5'h3 == out ? Qh_3_io_cmd_out_valid : _io_cmd_out_valid_T_5; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_9 = 5'h4 == out ? Qh_4_io_cmd_out_valid : _io_cmd_out_valid_T_7; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_11 = 5'h5 == out ? Qh_5_io_cmd_out_valid : _io_cmd_out_valid_T_9; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_13 = 5'h6 == out ? Qh_6_io_cmd_out_valid : _io_cmd_out_valid_T_11; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_15 = 5'h7 == out ? Qh_7_io_cmd_out_valid : _io_cmd_out_valid_T_13; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_17 = 5'h8 == out ? Qh_8_io_cmd_out_valid : _io_cmd_out_valid_T_15; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_19 = 5'h9 == out ? Qh_9_io_cmd_out_valid : _io_cmd_out_valid_T_17; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_21 = 5'ha == out ? Qh_10_io_cmd_out_valid : _io_cmd_out_valid_T_19; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_23 = 5'hb == out ? Qh_11_io_cmd_out_valid : _io_cmd_out_valid_T_21; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_25 = 5'hc == out ? Qh_12_io_cmd_out_valid : _io_cmd_out_valid_T_23; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_27 = 5'hd == out ? Qh_13_io_cmd_out_valid : _io_cmd_out_valid_T_25; // @[Mux.scala 80:57]
  wire  _io_cmd_out_valid_T_29 = 5'he == out ? Qh_14_io_cmd_out_valid : _io_cmd_out_valid_T_27; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_1 = Qh_0_io_c2h_length; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_3 = 5'h1 == out ? Qh_1_io_c2h_length : _io_c2h_length_T_1; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_5 = 5'h2 == out ? Qh_2_io_c2h_length : _io_c2h_length_T_3; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_7 = 5'h3 == out ? Qh_3_io_c2h_length : _io_c2h_length_T_5; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_9 = 5'h4 == out ? Qh_4_io_c2h_length : _io_c2h_length_T_7; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_11 = 5'h5 == out ? Qh_5_io_c2h_length : _io_c2h_length_T_9; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_13 = 5'h6 == out ? Qh_6_io_c2h_length : _io_c2h_length_T_11; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_15 = 5'h7 == out ? Qh_7_io_c2h_length : _io_c2h_length_T_13; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_17 = 5'h8 == out ? Qh_8_io_c2h_length : _io_c2h_length_T_15; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_19 = 5'h9 == out ? Qh_9_io_c2h_length : _io_c2h_length_T_17; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_21 = 5'ha == out ? Qh_10_io_c2h_length : _io_c2h_length_T_19; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_23 = 5'hb == out ? Qh_11_io_c2h_length : _io_c2h_length_T_21; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_25 = 5'hc == out ? Qh_12_io_c2h_length : _io_c2h_length_T_23; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_27 = 5'hd == out ? Qh_13_io_c2h_length : _io_c2h_length_T_25; // @[Mux.scala 80:57]
  wire [31:0] _io_c2h_length_T_29 = 5'he == out ? Qh_14_io_c2h_length : _io_c2h_length_T_27; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_3 = 5'h1 == out ? Qh_1_io_m2h_complete : Qh_0_io_m2h_complete; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_5 = 5'h2 == out ? Qh_2_io_m2h_complete : _io_m2h_complete_T_3; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_7 = 5'h3 == out ? Qh_3_io_m2h_complete : _io_m2h_complete_T_5; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_9 = 5'h4 == out ? Qh_4_io_m2h_complete : _io_m2h_complete_T_7; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_11 = 5'h5 == out ? Qh_5_io_m2h_complete : _io_m2h_complete_T_9; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_13 = 5'h6 == out ? Qh_6_io_m2h_complete : _io_m2h_complete_T_11; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_15 = 5'h7 == out ? Qh_7_io_m2h_complete : _io_m2h_complete_T_13; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_17 = 5'h8 == out ? Qh_8_io_m2h_complete : _io_m2h_complete_T_15; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_19 = 5'h9 == out ? Qh_9_io_m2h_complete : _io_m2h_complete_T_17; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_21 = 5'ha == out ? Qh_10_io_m2h_complete : _io_m2h_complete_T_19; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_23 = 5'hb == out ? Qh_11_io_m2h_complete : _io_m2h_complete_T_21; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_25 = 5'hc == out ? Qh_12_io_m2h_complete : _io_m2h_complete_T_23; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_27 = 5'hd == out ? Qh_13_io_m2h_complete : _io_m2h_complete_T_25; // @[Mux.scala 80:57]
  wire  _io_m2h_complete_T_29 = 5'he == out ? Qh_14_io_m2h_complete : _io_m2h_complete_T_27; // @[Mux.scala 80:57]
  wire  _io_last_T_3 = 5'h1 == out ? Qh_1_io_last : Qh_0_io_last; // @[Mux.scala 80:57]
  wire  _io_last_T_5 = 5'h2 == out ? Qh_2_io_last : _io_last_T_3; // @[Mux.scala 80:57]
  wire  _io_last_T_7 = 5'h3 == out ? Qh_3_io_last : _io_last_T_5; // @[Mux.scala 80:57]
  wire  _io_last_T_9 = 5'h4 == out ? Qh_4_io_last : _io_last_T_7; // @[Mux.scala 80:57]
  wire  _io_last_T_11 = 5'h5 == out ? Qh_5_io_last : _io_last_T_9; // @[Mux.scala 80:57]
  wire  _io_last_T_13 = 5'h6 == out ? Qh_6_io_last : _io_last_T_11; // @[Mux.scala 80:57]
  wire  _io_last_T_15 = 5'h7 == out ? Qh_7_io_last : _io_last_T_13; // @[Mux.scala 80:57]
  wire  _io_last_T_17 = 5'h8 == out ? Qh_8_io_last : _io_last_T_15; // @[Mux.scala 80:57]
  wire  _io_last_T_19 = 5'h9 == out ? Qh_9_io_last : _io_last_T_17; // @[Mux.scala 80:57]
  wire  _io_last_T_21 = 5'ha == out ? Qh_10_io_last : _io_last_T_19; // @[Mux.scala 80:57]
  wire  _io_last_T_23 = 5'hb == out ? Qh_11_io_last : _io_last_T_21; // @[Mux.scala 80:57]
  wire  _io_last_T_25 = 5'hc == out ? Qh_12_io_last : _io_last_T_23; // @[Mux.scala 80:57]
  wire  _io_last_T_27 = 5'hd == out ? Qh_13_io_last : _io_last_T_25; // @[Mux.scala 80:57]
  wire  _io_last_T_29 = 5'he == out ? Qh_14_io_last : _io_last_T_27; // @[Mux.scala 80:57]
  XQueue_18 Q_0 ( // @[XQueue.scala 35:23]
    .clock(Q_0_clock),
    .reset(Q_0_reset),
    .io_in_valid(Q_0_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_0_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_0_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_0_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_0_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_0_io_in_bits_pkt_size),
    .io_out_ready(Q_0_io_out_ready),
    .io_out_valid(Q_0_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_0_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_0_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_0_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_0_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_0_io_out_bits_pkt_size)
  );
  XQueue_18 Q_1 ( // @[XQueue.scala 35:23]
    .clock(Q_1_clock),
    .reset(Q_1_reset),
    .io_in_valid(Q_1_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_1_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_1_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_1_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_1_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_1_io_in_bits_pkt_size),
    .io_out_ready(Q_1_io_out_ready),
    .io_out_valid(Q_1_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_1_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_1_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_1_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_1_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_1_io_out_bits_pkt_size)
  );
  XQueue_18 Q_2 ( // @[XQueue.scala 35:23]
    .clock(Q_2_clock),
    .reset(Q_2_reset),
    .io_in_valid(Q_2_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_2_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_2_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_2_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_2_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_2_io_in_bits_pkt_size),
    .io_out_ready(Q_2_io_out_ready),
    .io_out_valid(Q_2_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_2_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_2_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_2_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_2_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_2_io_out_bits_pkt_size)
  );
  XQueue_18 Q_3 ( // @[XQueue.scala 35:23]
    .clock(Q_3_clock),
    .reset(Q_3_reset),
    .io_in_valid(Q_3_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_3_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_3_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_3_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_3_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_3_io_in_bits_pkt_size),
    .io_out_ready(Q_3_io_out_ready),
    .io_out_valid(Q_3_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_3_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_3_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_3_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_3_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_3_io_out_bits_pkt_size)
  );
  XQueue_18 Q_4 ( // @[XQueue.scala 35:23]
    .clock(Q_4_clock),
    .reset(Q_4_reset),
    .io_in_valid(Q_4_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_4_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_4_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_4_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_4_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_4_io_in_bits_pkt_size),
    .io_out_ready(Q_4_io_out_ready),
    .io_out_valid(Q_4_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_4_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_4_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_4_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_4_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_4_io_out_bits_pkt_size)
  );
  XQueue_18 Q_5 ( // @[XQueue.scala 35:23]
    .clock(Q_5_clock),
    .reset(Q_5_reset),
    .io_in_valid(Q_5_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_5_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_5_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_5_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_5_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_5_io_in_bits_pkt_size),
    .io_out_ready(Q_5_io_out_ready),
    .io_out_valid(Q_5_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_5_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_5_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_5_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_5_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_5_io_out_bits_pkt_size)
  );
  XQueue_18 Q_6 ( // @[XQueue.scala 35:23]
    .clock(Q_6_clock),
    .reset(Q_6_reset),
    .io_in_valid(Q_6_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_6_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_6_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_6_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_6_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_6_io_in_bits_pkt_size),
    .io_out_ready(Q_6_io_out_ready),
    .io_out_valid(Q_6_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_6_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_6_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_6_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_6_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_6_io_out_bits_pkt_size)
  );
  XQueue_18 Q_7 ( // @[XQueue.scala 35:23]
    .clock(Q_7_clock),
    .reset(Q_7_reset),
    .io_in_valid(Q_7_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_7_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_7_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_7_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_7_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_7_io_in_bits_pkt_size),
    .io_out_ready(Q_7_io_out_ready),
    .io_out_valid(Q_7_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_7_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_7_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_7_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_7_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_7_io_out_bits_pkt_size)
  );
  XQueue_18 Q_8 ( // @[XQueue.scala 35:23]
    .clock(Q_8_clock),
    .reset(Q_8_reset),
    .io_in_valid(Q_8_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_8_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_8_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_8_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_8_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_8_io_in_bits_pkt_size),
    .io_out_ready(Q_8_io_out_ready),
    .io_out_valid(Q_8_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_8_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_8_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_8_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_8_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_8_io_out_bits_pkt_size)
  );
  XQueue_18 Q_9 ( // @[XQueue.scala 35:23]
    .clock(Q_9_clock),
    .reset(Q_9_reset),
    .io_in_valid(Q_9_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_9_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_9_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_9_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_9_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_9_io_in_bits_pkt_size),
    .io_out_ready(Q_9_io_out_ready),
    .io_out_valid(Q_9_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_9_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_9_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_9_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_9_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_9_io_out_bits_pkt_size)
  );
  XQueue_18 Q_10 ( // @[XQueue.scala 35:23]
    .clock(Q_10_clock),
    .reset(Q_10_reset),
    .io_in_valid(Q_10_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_10_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_10_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_10_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_10_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_10_io_in_bits_pkt_size),
    .io_out_ready(Q_10_io_out_ready),
    .io_out_valid(Q_10_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_10_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_10_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_10_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_10_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_10_io_out_bits_pkt_size)
  );
  XQueue_18 Q_11 ( // @[XQueue.scala 35:23]
    .clock(Q_11_clock),
    .reset(Q_11_reset),
    .io_in_valid(Q_11_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_11_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_11_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_11_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_11_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_11_io_in_bits_pkt_size),
    .io_out_ready(Q_11_io_out_ready),
    .io_out_valid(Q_11_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_11_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_11_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_11_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_11_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_11_io_out_bits_pkt_size)
  );
  XQueue_18 Q_12 ( // @[XQueue.scala 35:23]
    .clock(Q_12_clock),
    .reset(Q_12_reset),
    .io_in_valid(Q_12_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_12_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_12_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_12_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_12_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_12_io_in_bits_pkt_size),
    .io_out_ready(Q_12_io_out_ready),
    .io_out_valid(Q_12_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_12_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_12_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_12_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_12_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_12_io_out_bits_pkt_size)
  );
  XQueue_18 Q_13 ( // @[XQueue.scala 35:23]
    .clock(Q_13_clock),
    .reset(Q_13_reset),
    .io_in_valid(Q_13_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_13_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_13_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_13_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_13_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_13_io_in_bits_pkt_size),
    .io_out_ready(Q_13_io_out_ready),
    .io_out_valid(Q_13_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_13_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_13_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_13_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_13_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_13_io_out_bits_pkt_size)
  );
  XQueue_18 Q_14 ( // @[XQueue.scala 35:23]
    .clock(Q_14_clock),
    .reset(Q_14_reset),
    .io_in_valid(Q_14_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_14_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_14_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_14_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_14_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_14_io_in_bits_pkt_size),
    .io_out_ready(Q_14_io_out_ready),
    .io_out_valid(Q_14_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_14_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_14_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_14_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_14_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_14_io_out_bits_pkt_size)
  );
  XQueue_18 Q_15 ( // @[XQueue.scala 35:23]
    .clock(Q_15_clock),
    .reset(Q_15_reset),
    .io_in_valid(Q_15_io_in_valid),
    .io_in_bits_c2h_start_addr(Q_15_io_in_bits_c2h_start_addr),
    .io_in_bits_m2h_start_addr(Q_15_io_in_bits_m2h_start_addr),
    .io_in_bits_m2h_length(Q_15_io_in_bits_m2h_length),
    .io_in_bits_c2h_cpt_addr(Q_15_io_in_bits_c2h_cpt_addr),
    .io_in_bits_pkt_size(Q_15_io_in_bits_pkt_size),
    .io_out_ready(Q_15_io_out_ready),
    .io_out_valid(Q_15_io_out_valid),
    .io_out_bits_c2h_start_addr(Q_15_io_out_bits_c2h_start_addr),
    .io_out_bits_m2h_start_addr(Q_15_io_out_bits_m2h_start_addr),
    .io_out_bits_m2h_length(Q_15_io_out_bits_m2h_length),
    .io_out_bits_c2h_cpt_addr(Q_15_io_out_bits_c2h_cpt_addr),
    .io_out_bits_pkt_size(Q_15_io_out_bits_pkt_size)
  );
  d2hcmdqueuehead Qh_0 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_0_clock),
    .reset(Qh_0_reset),
    .io_cmd_in_ready(Qh_0_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_0_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_0_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_0_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_0_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_0_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_0_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_0_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_0_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_0_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_0_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_0_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_0_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_0_io_c2h_length),
    .io_m2h_complete(Qh_0_io_m2h_complete),
    .io_c2h_finish(Qh_0_io_c2h_finish),
    .io_m2h_finish(Qh_0_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_0_io_m2h_cpt_complete),
    .io_last(Qh_0_io_last),
    .io_working(Qh_0_io_working),
    .io_continue(Qh_0_io_continue)
  );
  d2hcmdqueuehead Qh_1 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_1_clock),
    .reset(Qh_1_reset),
    .io_cmd_in_ready(Qh_1_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_1_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_1_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_1_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_1_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_1_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_1_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_1_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_1_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_1_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_1_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_1_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_1_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_1_io_c2h_length),
    .io_m2h_complete(Qh_1_io_m2h_complete),
    .io_c2h_finish(Qh_1_io_c2h_finish),
    .io_m2h_finish(Qh_1_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_1_io_m2h_cpt_complete),
    .io_last(Qh_1_io_last),
    .io_working(Qh_1_io_working),
    .io_continue(Qh_1_io_continue)
  );
  d2hcmdqueuehead Qh_2 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_2_clock),
    .reset(Qh_2_reset),
    .io_cmd_in_ready(Qh_2_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_2_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_2_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_2_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_2_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_2_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_2_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_2_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_2_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_2_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_2_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_2_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_2_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_2_io_c2h_length),
    .io_m2h_complete(Qh_2_io_m2h_complete),
    .io_c2h_finish(Qh_2_io_c2h_finish),
    .io_m2h_finish(Qh_2_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_2_io_m2h_cpt_complete),
    .io_last(Qh_2_io_last),
    .io_working(Qh_2_io_working),
    .io_continue(Qh_2_io_continue)
  );
  d2hcmdqueuehead Qh_3 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_3_clock),
    .reset(Qh_3_reset),
    .io_cmd_in_ready(Qh_3_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_3_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_3_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_3_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_3_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_3_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_3_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_3_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_3_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_3_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_3_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_3_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_3_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_3_io_c2h_length),
    .io_m2h_complete(Qh_3_io_m2h_complete),
    .io_c2h_finish(Qh_3_io_c2h_finish),
    .io_m2h_finish(Qh_3_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_3_io_m2h_cpt_complete),
    .io_last(Qh_3_io_last),
    .io_working(Qh_3_io_working),
    .io_continue(Qh_3_io_continue)
  );
  d2hcmdqueuehead Qh_4 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_4_clock),
    .reset(Qh_4_reset),
    .io_cmd_in_ready(Qh_4_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_4_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_4_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_4_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_4_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_4_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_4_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_4_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_4_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_4_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_4_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_4_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_4_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_4_io_c2h_length),
    .io_m2h_complete(Qh_4_io_m2h_complete),
    .io_c2h_finish(Qh_4_io_c2h_finish),
    .io_m2h_finish(Qh_4_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_4_io_m2h_cpt_complete),
    .io_last(Qh_4_io_last),
    .io_working(Qh_4_io_working),
    .io_continue(Qh_4_io_continue)
  );
  d2hcmdqueuehead Qh_5 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_5_clock),
    .reset(Qh_5_reset),
    .io_cmd_in_ready(Qh_5_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_5_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_5_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_5_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_5_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_5_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_5_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_5_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_5_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_5_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_5_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_5_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_5_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_5_io_c2h_length),
    .io_m2h_complete(Qh_5_io_m2h_complete),
    .io_c2h_finish(Qh_5_io_c2h_finish),
    .io_m2h_finish(Qh_5_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_5_io_m2h_cpt_complete),
    .io_last(Qh_5_io_last),
    .io_working(Qh_5_io_working),
    .io_continue(Qh_5_io_continue)
  );
  d2hcmdqueuehead Qh_6 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_6_clock),
    .reset(Qh_6_reset),
    .io_cmd_in_ready(Qh_6_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_6_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_6_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_6_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_6_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_6_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_6_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_6_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_6_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_6_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_6_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_6_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_6_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_6_io_c2h_length),
    .io_m2h_complete(Qh_6_io_m2h_complete),
    .io_c2h_finish(Qh_6_io_c2h_finish),
    .io_m2h_finish(Qh_6_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_6_io_m2h_cpt_complete),
    .io_last(Qh_6_io_last),
    .io_working(Qh_6_io_working),
    .io_continue(Qh_6_io_continue)
  );
  d2hcmdqueuehead Qh_7 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_7_clock),
    .reset(Qh_7_reset),
    .io_cmd_in_ready(Qh_7_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_7_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_7_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_7_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_7_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_7_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_7_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_7_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_7_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_7_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_7_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_7_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_7_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_7_io_c2h_length),
    .io_m2h_complete(Qh_7_io_m2h_complete),
    .io_c2h_finish(Qh_7_io_c2h_finish),
    .io_m2h_finish(Qh_7_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_7_io_m2h_cpt_complete),
    .io_last(Qh_7_io_last),
    .io_working(Qh_7_io_working),
    .io_continue(Qh_7_io_continue)
  );
  d2hcmdqueuehead Qh_8 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_8_clock),
    .reset(Qh_8_reset),
    .io_cmd_in_ready(Qh_8_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_8_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_8_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_8_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_8_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_8_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_8_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_8_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_8_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_8_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_8_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_8_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_8_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_8_io_c2h_length),
    .io_m2h_complete(Qh_8_io_m2h_complete),
    .io_c2h_finish(Qh_8_io_c2h_finish),
    .io_m2h_finish(Qh_8_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_8_io_m2h_cpt_complete),
    .io_last(Qh_8_io_last),
    .io_working(Qh_8_io_working),
    .io_continue(Qh_8_io_continue)
  );
  d2hcmdqueuehead Qh_9 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_9_clock),
    .reset(Qh_9_reset),
    .io_cmd_in_ready(Qh_9_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_9_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_9_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_9_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_9_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_9_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_9_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_9_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_9_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_9_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_9_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_9_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_9_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_9_io_c2h_length),
    .io_m2h_complete(Qh_9_io_m2h_complete),
    .io_c2h_finish(Qh_9_io_c2h_finish),
    .io_m2h_finish(Qh_9_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_9_io_m2h_cpt_complete),
    .io_last(Qh_9_io_last),
    .io_working(Qh_9_io_working),
    .io_continue(Qh_9_io_continue)
  );
  d2hcmdqueuehead Qh_10 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_10_clock),
    .reset(Qh_10_reset),
    .io_cmd_in_ready(Qh_10_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_10_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_10_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_10_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_10_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_10_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_10_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_10_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_10_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_10_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_10_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_10_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_10_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_10_io_c2h_length),
    .io_m2h_complete(Qh_10_io_m2h_complete),
    .io_c2h_finish(Qh_10_io_c2h_finish),
    .io_m2h_finish(Qh_10_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_10_io_m2h_cpt_complete),
    .io_last(Qh_10_io_last),
    .io_working(Qh_10_io_working),
    .io_continue(Qh_10_io_continue)
  );
  d2hcmdqueuehead Qh_11 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_11_clock),
    .reset(Qh_11_reset),
    .io_cmd_in_ready(Qh_11_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_11_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_11_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_11_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_11_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_11_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_11_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_11_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_11_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_11_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_11_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_11_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_11_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_11_io_c2h_length),
    .io_m2h_complete(Qh_11_io_m2h_complete),
    .io_c2h_finish(Qh_11_io_c2h_finish),
    .io_m2h_finish(Qh_11_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_11_io_m2h_cpt_complete),
    .io_last(Qh_11_io_last),
    .io_working(Qh_11_io_working),
    .io_continue(Qh_11_io_continue)
  );
  d2hcmdqueuehead Qh_12 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_12_clock),
    .reset(Qh_12_reset),
    .io_cmd_in_ready(Qh_12_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_12_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_12_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_12_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_12_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_12_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_12_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_12_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_12_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_12_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_12_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_12_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_12_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_12_io_c2h_length),
    .io_m2h_complete(Qh_12_io_m2h_complete),
    .io_c2h_finish(Qh_12_io_c2h_finish),
    .io_m2h_finish(Qh_12_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_12_io_m2h_cpt_complete),
    .io_last(Qh_12_io_last),
    .io_working(Qh_12_io_working),
    .io_continue(Qh_12_io_continue)
  );
  d2hcmdqueuehead Qh_13 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_13_clock),
    .reset(Qh_13_reset),
    .io_cmd_in_ready(Qh_13_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_13_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_13_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_13_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_13_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_13_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_13_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_13_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_13_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_13_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_13_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_13_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_13_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_13_io_c2h_length),
    .io_m2h_complete(Qh_13_io_m2h_complete),
    .io_c2h_finish(Qh_13_io_c2h_finish),
    .io_m2h_finish(Qh_13_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_13_io_m2h_cpt_complete),
    .io_last(Qh_13_io_last),
    .io_working(Qh_13_io_working),
    .io_continue(Qh_13_io_continue)
  );
  d2hcmdqueuehead Qh_14 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_14_clock),
    .reset(Qh_14_reset),
    .io_cmd_in_ready(Qh_14_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_14_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_14_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_14_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_14_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_14_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_14_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_14_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_14_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_14_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_14_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_14_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_14_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_14_io_c2h_length),
    .io_m2h_complete(Qh_14_io_m2h_complete),
    .io_c2h_finish(Qh_14_io_c2h_finish),
    .io_m2h_finish(Qh_14_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_14_io_m2h_cpt_complete),
    .io_last(Qh_14_io_last),
    .io_working(Qh_14_io_working),
    .io_continue(Qh_14_io_continue)
  );
  d2hcmdqueuehead Qh_15 ( // @[d2hcmdqueue.scala 35:45]
    .clock(Qh_15_clock),
    .reset(Qh_15_reset),
    .io_cmd_in_ready(Qh_15_io_cmd_in_ready),
    .io_cmd_in_valid(Qh_15_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(Qh_15_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(Qh_15_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(Qh_15_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(Qh_15_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(Qh_15_io_cmd_in_bits_pkt_size),
    .io_cmd_out_ready(Qh_15_io_cmd_out_ready),
    .io_cmd_out_valid(Qh_15_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(Qh_15_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(Qh_15_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(Qh_15_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(Qh_15_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(Qh_15_io_c2h_length),
    .io_m2h_complete(Qh_15_io_m2h_complete),
    .io_c2h_finish(Qh_15_io_c2h_finish),
    .io_m2h_finish(Qh_15_io_m2h_finish),
    .io_m2h_cpt_complete(Qh_15_io_m2h_cpt_complete),
    .io_last(Qh_15_io_last),
    .io_working(Qh_15_io_working),
    .io_continue(Qh_15_io_continue)
  );
  assign io_cmd_out_valid = 5'hf == out ? Qh_15_io_cmd_out_valid : _io_cmd_out_valid_T_29; // @[Mux.scala 80:57]
  assign io_cmd_out_bits_c2h_start_addr = 5'hf == out ? Qh_15_io_cmd_out_bits_c2h_start_addr :
    _io_cmd_out_bits_T_29_c2h_start_addr; // @[Mux.scala 80:57]
  assign io_cmd_out_bits_m2h_start_addr = 5'hf == out ? Qh_15_io_cmd_out_bits_m2h_start_addr :
    _io_cmd_out_bits_T_29_m2h_start_addr; // @[Mux.scala 80:57]
  assign io_cmd_out_bits_m2h_length = 5'hf == out ? Qh_15_io_cmd_out_bits_m2h_length : _io_cmd_out_bits_T_29_m2h_length; // @[Mux.scala 80:57]
  assign io_cmd_out_bits_c2h_cpt_addr = 5'hf == out ? Qh_15_io_cmd_out_bits_c2h_cpt_addr :
    _io_cmd_out_bits_T_29_c2h_cpt_addr; // @[Mux.scala 80:57]
  assign io_c2h_length = 5'hf == out ? Qh_15_io_c2h_length : _io_c2h_length_T_29; // @[Mux.scala 80:57]
  assign io_m2h_complete = 5'hf == out ? Qh_15_io_m2h_complete : _io_m2h_complete_T_29; // @[Mux.scala 80:57]
  assign io_h2m_complete = h2m_complete; // @[d2hcmdqueue.scala 48:21]
  assign io_last = 5'hf == out ? Qh_15_io_last : _io_last_T_29; // @[Mux.scala 80:57]
  assign io_counter = counter; // @[d2hcmdqueue.scala 38:16]
  assign Q_0_clock = clock;
  assign Q_0_reset = reset;
  assign Q_0_io_in_valid = io_cmd_in_valid & io_qin[0]; // @[d2hcmdqueue.scala 60:56]
  assign Q_0_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_0_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_0_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_0_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_0_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_0_io_out_ready = Qh_0_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_1_clock = clock;
  assign Q_1_reset = reset;
  assign Q_1_io_in_valid = io_cmd_in_valid & io_qin[1]; // @[d2hcmdqueue.scala 60:56]
  assign Q_1_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_1_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_1_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_1_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_1_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_1_io_out_ready = Qh_1_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_2_clock = clock;
  assign Q_2_reset = reset;
  assign Q_2_io_in_valid = io_cmd_in_valid & io_qin[2]; // @[d2hcmdqueue.scala 60:56]
  assign Q_2_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_2_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_2_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_2_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_2_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_2_io_out_ready = Qh_2_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_3_clock = clock;
  assign Q_3_reset = reset;
  assign Q_3_io_in_valid = io_cmd_in_valid & io_qin[3]; // @[d2hcmdqueue.scala 60:56]
  assign Q_3_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_3_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_3_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_3_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_3_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_3_io_out_ready = Qh_3_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_4_clock = clock;
  assign Q_4_reset = reset;
  assign Q_4_io_in_valid = io_cmd_in_valid & io_qin[4]; // @[d2hcmdqueue.scala 60:56]
  assign Q_4_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_4_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_4_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_4_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_4_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_4_io_out_ready = Qh_4_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_5_clock = clock;
  assign Q_5_reset = reset;
  assign Q_5_io_in_valid = io_cmd_in_valid & io_qin[5]; // @[d2hcmdqueue.scala 60:56]
  assign Q_5_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_5_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_5_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_5_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_5_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_5_io_out_ready = Qh_5_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_6_clock = clock;
  assign Q_6_reset = reset;
  assign Q_6_io_in_valid = io_cmd_in_valid & io_qin[6]; // @[d2hcmdqueue.scala 60:56]
  assign Q_6_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_6_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_6_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_6_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_6_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_6_io_out_ready = Qh_6_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_7_clock = clock;
  assign Q_7_reset = reset;
  assign Q_7_io_in_valid = io_cmd_in_valid & io_qin[7]; // @[d2hcmdqueue.scala 60:56]
  assign Q_7_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_7_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_7_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_7_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_7_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_7_io_out_ready = Qh_7_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_8_clock = clock;
  assign Q_8_reset = reset;
  assign Q_8_io_in_valid = io_cmd_in_valid & io_qin[8]; // @[d2hcmdqueue.scala 60:56]
  assign Q_8_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_8_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_8_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_8_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_8_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_8_io_out_ready = Qh_8_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_9_clock = clock;
  assign Q_9_reset = reset;
  assign Q_9_io_in_valid = io_cmd_in_valid & io_qin[9]; // @[d2hcmdqueue.scala 60:56]
  assign Q_9_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_9_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_9_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_9_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_9_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_9_io_out_ready = Qh_9_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_10_clock = clock;
  assign Q_10_reset = reset;
  assign Q_10_io_in_valid = io_cmd_in_valid & io_qin[10]; // @[d2hcmdqueue.scala 60:56]
  assign Q_10_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_10_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_10_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_10_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_10_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_10_io_out_ready = Qh_10_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_11_clock = clock;
  assign Q_11_reset = reset;
  assign Q_11_io_in_valid = io_cmd_in_valid & io_qin[11]; // @[d2hcmdqueue.scala 60:56]
  assign Q_11_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_11_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_11_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_11_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_11_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_11_io_out_ready = Qh_11_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_12_clock = clock;
  assign Q_12_reset = reset;
  assign Q_12_io_in_valid = io_cmd_in_valid & io_qin[12]; // @[d2hcmdqueue.scala 60:56]
  assign Q_12_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_12_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_12_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_12_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_12_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_12_io_out_ready = Qh_12_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_13_clock = clock;
  assign Q_13_reset = reset;
  assign Q_13_io_in_valid = io_cmd_in_valid & io_qin[13]; // @[d2hcmdqueue.scala 60:56]
  assign Q_13_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_13_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_13_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_13_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_13_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_13_io_out_ready = Qh_13_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_14_clock = clock;
  assign Q_14_reset = reset;
  assign Q_14_io_in_valid = io_cmd_in_valid & io_qin[14]; // @[d2hcmdqueue.scala 60:56]
  assign Q_14_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_14_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_14_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_14_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_14_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_14_io_out_ready = Qh_14_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Q_15_clock = clock;
  assign Q_15_reset = reset;
  assign Q_15_io_in_valid = io_cmd_in_valid & io_qin[15]; // @[d2hcmdqueue.scala 60:56]
  assign Q_15_io_in_bits_c2h_start_addr = io_cmd_in_bits_c2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_15_io_in_bits_m2h_start_addr = io_cmd_in_bits_m2h_start_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_15_io_in_bits_m2h_length = io_cmd_in_bits_m2h_length; // @[d2hcmdqueue.scala 61:37]
  assign Q_15_io_in_bits_c2h_cpt_addr = io_cmd_in_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 61:37]
  assign Q_15_io_in_bits_pkt_size = io_cmd_in_bits_pkt_size; // @[d2hcmdqueue.scala 61:37]
  assign Q_15_io_out_ready = Qh_15_io_cmd_in_ready; // @[d2hcmdqueue.scala 62:37]
  assign Qh_0_clock = clock;
  assign Qh_0_reset = reset;
  assign Qh_0_io_cmd_in_valid = Q_0_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_0_io_cmd_in_bits_c2h_start_addr = Q_0_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_0_io_cmd_in_bits_m2h_start_addr = Q_0_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_0_io_cmd_in_bits_m2h_length = Q_0_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_0_io_cmd_in_bits_c2h_cpt_addr = Q_0_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_0_io_cmd_in_bits_pkt_size = Q_0_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_0_io_cmd_out_ready = io_cmd_out_ready & out == 5'h0; // @[d2hcmdqueue.scala 63:57]
  assign Qh_0_io_c2h_finish = io_c2h_finish & _Qh_0_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_0_io_m2h_finish = io_m2h_finish & _Qh_0_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_0_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_0_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_1_clock = clock;
  assign Qh_1_reset = reset;
  assign Qh_1_io_cmd_in_valid = Q_1_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_1_io_cmd_in_bits_c2h_start_addr = Q_1_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_1_io_cmd_in_bits_m2h_start_addr = Q_1_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_1_io_cmd_in_bits_m2h_length = Q_1_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_1_io_cmd_in_bits_c2h_cpt_addr = Q_1_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_1_io_cmd_in_bits_pkt_size = Q_1_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_1_io_cmd_out_ready = io_cmd_out_ready & out == 5'h1; // @[d2hcmdqueue.scala 63:57]
  assign Qh_1_io_c2h_finish = io_c2h_finish & _Qh_1_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_1_io_m2h_finish = io_m2h_finish & _Qh_1_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_1_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_1_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_2_clock = clock;
  assign Qh_2_reset = reset;
  assign Qh_2_io_cmd_in_valid = Q_2_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_2_io_cmd_in_bits_c2h_start_addr = Q_2_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_2_io_cmd_in_bits_m2h_start_addr = Q_2_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_2_io_cmd_in_bits_m2h_length = Q_2_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_2_io_cmd_in_bits_c2h_cpt_addr = Q_2_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_2_io_cmd_in_bits_pkt_size = Q_2_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_2_io_cmd_out_ready = io_cmd_out_ready & out == 5'h2; // @[d2hcmdqueue.scala 63:57]
  assign Qh_2_io_c2h_finish = io_c2h_finish & _Qh_2_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_2_io_m2h_finish = io_m2h_finish & _Qh_2_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_2_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_2_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_3_clock = clock;
  assign Qh_3_reset = reset;
  assign Qh_3_io_cmd_in_valid = Q_3_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_3_io_cmd_in_bits_c2h_start_addr = Q_3_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_3_io_cmd_in_bits_m2h_start_addr = Q_3_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_3_io_cmd_in_bits_m2h_length = Q_3_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_3_io_cmd_in_bits_c2h_cpt_addr = Q_3_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_3_io_cmd_in_bits_pkt_size = Q_3_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_3_io_cmd_out_ready = io_cmd_out_ready & out == 5'h3; // @[d2hcmdqueue.scala 63:57]
  assign Qh_3_io_c2h_finish = io_c2h_finish & _Qh_3_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_3_io_m2h_finish = io_m2h_finish & _Qh_3_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_3_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_3_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_4_clock = clock;
  assign Qh_4_reset = reset;
  assign Qh_4_io_cmd_in_valid = Q_4_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_4_io_cmd_in_bits_c2h_start_addr = Q_4_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_4_io_cmd_in_bits_m2h_start_addr = Q_4_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_4_io_cmd_in_bits_m2h_length = Q_4_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_4_io_cmd_in_bits_c2h_cpt_addr = Q_4_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_4_io_cmd_in_bits_pkt_size = Q_4_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_4_io_cmd_out_ready = io_cmd_out_ready & out == 5'h4; // @[d2hcmdqueue.scala 63:57]
  assign Qh_4_io_c2h_finish = io_c2h_finish & _Qh_4_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_4_io_m2h_finish = io_m2h_finish & _Qh_4_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_4_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_4_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_5_clock = clock;
  assign Qh_5_reset = reset;
  assign Qh_5_io_cmd_in_valid = Q_5_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_5_io_cmd_in_bits_c2h_start_addr = Q_5_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_5_io_cmd_in_bits_m2h_start_addr = Q_5_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_5_io_cmd_in_bits_m2h_length = Q_5_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_5_io_cmd_in_bits_c2h_cpt_addr = Q_5_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_5_io_cmd_in_bits_pkt_size = Q_5_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_5_io_cmd_out_ready = io_cmd_out_ready & out == 5'h5; // @[d2hcmdqueue.scala 63:57]
  assign Qh_5_io_c2h_finish = io_c2h_finish & _Qh_5_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_5_io_m2h_finish = io_m2h_finish & _Qh_5_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_5_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_5_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_6_clock = clock;
  assign Qh_6_reset = reset;
  assign Qh_6_io_cmd_in_valid = Q_6_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_6_io_cmd_in_bits_c2h_start_addr = Q_6_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_6_io_cmd_in_bits_m2h_start_addr = Q_6_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_6_io_cmd_in_bits_m2h_length = Q_6_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_6_io_cmd_in_bits_c2h_cpt_addr = Q_6_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_6_io_cmd_in_bits_pkt_size = Q_6_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_6_io_cmd_out_ready = io_cmd_out_ready & out == 5'h6; // @[d2hcmdqueue.scala 63:57]
  assign Qh_6_io_c2h_finish = io_c2h_finish & _Qh_6_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_6_io_m2h_finish = io_m2h_finish & _Qh_6_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_6_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_6_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_7_clock = clock;
  assign Qh_7_reset = reset;
  assign Qh_7_io_cmd_in_valid = Q_7_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_7_io_cmd_in_bits_c2h_start_addr = Q_7_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_7_io_cmd_in_bits_m2h_start_addr = Q_7_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_7_io_cmd_in_bits_m2h_length = Q_7_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_7_io_cmd_in_bits_c2h_cpt_addr = Q_7_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_7_io_cmd_in_bits_pkt_size = Q_7_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_7_io_cmd_out_ready = io_cmd_out_ready & out == 5'h7; // @[d2hcmdqueue.scala 63:57]
  assign Qh_7_io_c2h_finish = io_c2h_finish & _Qh_7_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_7_io_m2h_finish = io_m2h_finish & _Qh_7_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_7_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_7_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_8_clock = clock;
  assign Qh_8_reset = reset;
  assign Qh_8_io_cmd_in_valid = Q_8_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_8_io_cmd_in_bits_c2h_start_addr = Q_8_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_8_io_cmd_in_bits_m2h_start_addr = Q_8_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_8_io_cmd_in_bits_m2h_length = Q_8_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_8_io_cmd_in_bits_c2h_cpt_addr = Q_8_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_8_io_cmd_in_bits_pkt_size = Q_8_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_8_io_cmd_out_ready = io_cmd_out_ready & out == 5'h8; // @[d2hcmdqueue.scala 63:57]
  assign Qh_8_io_c2h_finish = io_c2h_finish & _Qh_8_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_8_io_m2h_finish = io_m2h_finish & _Qh_8_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_8_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_8_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_9_clock = clock;
  assign Qh_9_reset = reset;
  assign Qh_9_io_cmd_in_valid = Q_9_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_9_io_cmd_in_bits_c2h_start_addr = Q_9_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_9_io_cmd_in_bits_m2h_start_addr = Q_9_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_9_io_cmd_in_bits_m2h_length = Q_9_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_9_io_cmd_in_bits_c2h_cpt_addr = Q_9_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_9_io_cmd_in_bits_pkt_size = Q_9_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_9_io_cmd_out_ready = io_cmd_out_ready & out == 5'h9; // @[d2hcmdqueue.scala 63:57]
  assign Qh_9_io_c2h_finish = io_c2h_finish & _Qh_9_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_9_io_m2h_finish = io_m2h_finish & _Qh_9_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_9_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_9_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_10_clock = clock;
  assign Qh_10_reset = reset;
  assign Qh_10_io_cmd_in_valid = Q_10_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_10_io_cmd_in_bits_c2h_start_addr = Q_10_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_10_io_cmd_in_bits_m2h_start_addr = Q_10_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_10_io_cmd_in_bits_m2h_length = Q_10_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_10_io_cmd_in_bits_c2h_cpt_addr = Q_10_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_10_io_cmd_in_bits_pkt_size = Q_10_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_10_io_cmd_out_ready = io_cmd_out_ready & out == 5'ha; // @[d2hcmdqueue.scala 63:57]
  assign Qh_10_io_c2h_finish = io_c2h_finish & _Qh_10_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_10_io_m2h_finish = io_m2h_finish & _Qh_10_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_10_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_10_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_11_clock = clock;
  assign Qh_11_reset = reset;
  assign Qh_11_io_cmd_in_valid = Q_11_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_11_io_cmd_in_bits_c2h_start_addr = Q_11_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_11_io_cmd_in_bits_m2h_start_addr = Q_11_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_11_io_cmd_in_bits_m2h_length = Q_11_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_11_io_cmd_in_bits_c2h_cpt_addr = Q_11_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_11_io_cmd_in_bits_pkt_size = Q_11_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_11_io_cmd_out_ready = io_cmd_out_ready & out == 5'hb; // @[d2hcmdqueue.scala 63:57]
  assign Qh_11_io_c2h_finish = io_c2h_finish & _Qh_11_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_11_io_m2h_finish = io_m2h_finish & _Qh_11_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_11_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_11_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_12_clock = clock;
  assign Qh_12_reset = reset;
  assign Qh_12_io_cmd_in_valid = Q_12_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_12_io_cmd_in_bits_c2h_start_addr = Q_12_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_12_io_cmd_in_bits_m2h_start_addr = Q_12_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_12_io_cmd_in_bits_m2h_length = Q_12_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_12_io_cmd_in_bits_c2h_cpt_addr = Q_12_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_12_io_cmd_in_bits_pkt_size = Q_12_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_12_io_cmd_out_ready = io_cmd_out_ready & out == 5'hc; // @[d2hcmdqueue.scala 63:57]
  assign Qh_12_io_c2h_finish = io_c2h_finish & _Qh_12_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_12_io_m2h_finish = io_m2h_finish & _Qh_12_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_12_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_12_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_13_clock = clock;
  assign Qh_13_reset = reset;
  assign Qh_13_io_cmd_in_valid = Q_13_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_13_io_cmd_in_bits_c2h_start_addr = Q_13_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_13_io_cmd_in_bits_m2h_start_addr = Q_13_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_13_io_cmd_in_bits_m2h_length = Q_13_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_13_io_cmd_in_bits_c2h_cpt_addr = Q_13_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_13_io_cmd_in_bits_pkt_size = Q_13_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_13_io_cmd_out_ready = io_cmd_out_ready & out == 5'hd; // @[d2hcmdqueue.scala 63:57]
  assign Qh_13_io_c2h_finish = io_c2h_finish & _Qh_13_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_13_io_m2h_finish = io_m2h_finish & _Qh_13_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_13_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_13_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_14_clock = clock;
  assign Qh_14_reset = reset;
  assign Qh_14_io_cmd_in_valid = Q_14_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_14_io_cmd_in_bits_c2h_start_addr = Q_14_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_14_io_cmd_in_bits_m2h_start_addr = Q_14_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_14_io_cmd_in_bits_m2h_length = Q_14_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_14_io_cmd_in_bits_c2h_cpt_addr = Q_14_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_14_io_cmd_in_bits_pkt_size = Q_14_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_14_io_cmd_out_ready = io_cmd_out_ready & out == 5'he; // @[d2hcmdqueue.scala 63:57]
  assign Qh_14_io_c2h_finish = io_c2h_finish & _Qh_14_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_14_io_m2h_finish = io_m2h_finish & _Qh_14_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_14_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_14_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  assign Qh_15_clock = clock;
  assign Qh_15_reset = reset;
  assign Qh_15_io_cmd_in_valid = Q_15_io_out_valid; // @[d2hcmdqueue.scala 62:37]
  assign Qh_15_io_cmd_in_bits_c2h_start_addr = Q_15_io_out_bits_c2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_15_io_cmd_in_bits_m2h_start_addr = Q_15_io_out_bits_m2h_start_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_15_io_cmd_in_bits_m2h_length = Q_15_io_out_bits_m2h_length; // @[d2hcmdqueue.scala 62:37]
  assign Qh_15_io_cmd_in_bits_c2h_cpt_addr = Q_15_io_out_bits_c2h_cpt_addr; // @[d2hcmdqueue.scala 62:37]
  assign Qh_15_io_cmd_in_bits_pkt_size = Q_15_io_out_bits_pkt_size; // @[d2hcmdqueue.scala 62:37]
  assign Qh_15_io_cmd_out_ready = io_cmd_out_ready & out == 5'hf; // @[d2hcmdqueue.scala 63:57]
  assign Qh_15_io_c2h_finish = io_c2h_finish & _Qh_15_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 64:54]
  assign Qh_15_io_m2h_finish = io_m2h_finish & _Qh_15_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 65:54]
  assign Qh_15_io_m2h_cpt_complete = io_m2h_cpt_complete & _Qh_15_io_cmd_out_ready_T; // @[d2hcmdqueue.scala 66:60]
  always @(posedge clock) begin
    if (reset) begin // @[d2hcmdqueue.scala 37:26]
      counter <= 32'h0; // @[d2hcmdqueue.scala 37:26]
    end else if (_T) begin // @[d2hcmdqueue.scala 40:5]
      counter <= _counter_T_1; // @[d2hcmdqueue.scala 41:17]
    end
    if (reset) begin // @[d2hcmdqueue.scala 46:34]
      h2m_cpt_working <= 1'h0; // @[d2hcmdqueue.scala 46:34]
    end else if (out == 5'h1f) begin // @[d2hcmdqueue.scala 97:24]
      if (_T_441) begin // @[d2hcmdqueue.scala 107:13]
        h2m_cpt_working <= 1'h0; // @[d2hcmdqueue.scala 109:33]
      end else begin
        h2m_cpt_working <= _GEN_1;
      end
    end else begin
      h2m_cpt_working <= _GEN_1;
    end
    if (reset) begin // @[d2hcmdqueue.scala 47:31]
      h2m_complete <= 1'h0; // @[d2hcmdqueue.scala 47:31]
    end else if (out == 5'h1f) begin // @[d2hcmdqueue.scala 97:24]
      if (_T_441) begin // @[d2hcmdqueue.scala 107:13]
        h2m_complete <= 1'h0; // @[d2hcmdqueue.scala 108:30]
      end else if (!(_T_434)) begin // @[d2hcmdqueue.scala 99:13]
        h2m_complete <= _GEN_132;
      end
    end
    if (reset) begin // @[d2hcmdqueue.scala 54:23]
      out <= 5'h0; // @[d2hcmdqueue.scala 54:23]
    end else if (out == 5'h1f) begin // @[d2hcmdqueue.scala 97:24]
      if (_T_441) begin // @[d2hcmdqueue.scala 107:13]
        out <= next; // @[d2hcmdqueue.scala 110:21]
      end else begin
        out <= _GEN_126;
      end
    end else begin
      out <= _GEN_126;
    end
    if (reset) begin // @[d2hcmdqueue.scala 55:23]
      next <= 5'h0; // @[d2hcmdqueue.scala 55:23]
    end else if (_T_406 & next == 5'hf) begin // @[d2hcmdqueue.scala 89:58]
      next <= _GEN_4;
    end else if (Qh_15_io_continue & _Qh_15_io_cmd_out_ready_T & _T_4) begin // @[d2hcmdqueue.scala 78:77]
      next <= _GEN_4;
    end else if (_T_379 & next == 5'he) begin // @[d2hcmdqueue.scala 89:58]
      next <= _GEN_4;
    end else begin
      next <= _GEN_119;
    end
    if (reset) begin // @[d2hcmdqueue.scala 56:24]
      hold1 <= 5'h3; // @[d2hcmdqueue.scala 56:24]
    end else if (out == 5'h1f) begin // @[d2hcmdqueue.scala 97:24]
      if (_T_441) begin // @[d2hcmdqueue.scala 107:13]
        hold1 <= 5'h3; // @[d2hcmdqueue.scala 111:23]
      end else if (_T_434) begin // @[d2hcmdqueue.scala 99:13]
        hold1 <= _hold1_T_1; // @[d2hcmdqueue.scala 99:20]
      end
    end
    if (reset) begin // @[d2hcmdqueue.scala 57:24]
      hold2 <= 5'h3; // @[d2hcmdqueue.scala 57:24]
    end else if (out == 5'h1f) begin // @[d2hcmdqueue.scala 97:24]
      if (_T_441) begin // @[d2hcmdqueue.scala 107:13]
        hold2 <= 5'h3; // @[d2hcmdqueue.scala 112:23]
      end else if (!(_T_434)) begin // @[d2hcmdqueue.scala 99:13]
        hold2 <= _GEN_131;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  h2m_cpt_working = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  h2m_complete = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  out = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  next = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  hold1 = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  hold2 = _RAND_6[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module C2H(
  input         clock,
  input         reset,
  input  [63:0] io_start_addr,
  input  [31:0] io_length,
  input         io_start,
  input         io_c2h_cmd_ready,
  output        io_c2h_cmd_valid,
  output [63:0] io_c2h_cmd_bits_addr,
  output [6:0]  io_c2h_cmd_bits_pfch_tag,
  output [31:0] io_c2h_cmd_bits_len,
  input  [31:0] io_pfch_tag,
  output        io_complete,
  output [31:0] io_count_time,
  output [31:0] io_send_cmd_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] addr; // @[C2H.scala 23:50]
  reg [31:0] length; // @[C2H.scala 24:50]
  reg  valid_cmd; // @[C2H.scala 25:42]
  reg [31:0] count_time; // @[C2H.scala 29:42]
  reg [31:0] send_cmd_count; // @[C2H.scala 30:42]
  reg  complete; // @[C2H.scala 33:42]
  reg [3:0] hold; // @[C2H.scala 35:50]
  reg [1:0] state_cmd; // @[C2H.scala 48:42]
  wire  _T = 2'h0 == state_cmd; // @[Conditional.scala 37:30]
  wire  _GEN_1 = io_start ? 1'h0 : complete; // @[C2H.scala 53:39 C2H.scala 55:65 C2H.scala 33:42]
  wire  _T_1 = 2'h1 == state_cmd; // @[Conditional.scala 37:30]
  wire [31:0] _count_time_T_1 = count_time + 32'h1; // @[C2H.scala 64:79]
  wire  _T_2 = io_c2h_cmd_ready & io_c2h_cmd_valid; // @[Decoupled.scala 40:37]
  wire  _T_3 = 2'h2 == state_cmd; // @[Conditional.scala 37:30]
  wire [3:0] _hold_T_1 = hold - 4'h1; // @[C2H.scala 73:38]
  wire  _GEN_10 = hold == 4'h0 | complete; // @[C2H.scala 74:44 C2H.scala 75:65 C2H.scala 33:42]
  wire [1:0] _GEN_11 = hold == 4'h0 ? 2'h0 : state_cmd; // @[C2H.scala 74:44 C2H.scala 76:65 C2H.scala 48:42]
  wire  _GEN_13 = _T_3 ? _GEN_10 : complete; // @[Conditional.scala 39:67 C2H.scala 33:42]
  wire  _GEN_19 = _T_1 ? complete : _GEN_13; // @[Conditional.scala 39:67 C2H.scala 33:42]
  wire  _GEN_21 = _T ? _GEN_1 : _GEN_19; // @[Conditional.scala 40:58]
  wire [31:0] _send_cmd_count_T_1 = send_cmd_count + 32'h1; // @[C2H.scala 82:51]
  assign io_c2h_cmd_valid = valid_cmd; // @[C2H.scala 44:33]
  assign io_c2h_cmd_bits_addr = addr; // @[C2H.scala 41:33]
  assign io_c2h_cmd_bits_pfch_tag = io_pfch_tag[6:0]; // @[C2H.scala 42:33]
  assign io_c2h_cmd_bits_len = length; // @[C2H.scala 43:33]
  assign io_complete = complete; // @[C2H.scala 85:33]
  assign io_count_time = count_time; // @[C2H.scala 86:33]
  assign io_send_cmd_count = send_cmd_count; // @[C2H.scala 87:33]
  always @(posedge clock) begin
    if (reset) begin // @[C2H.scala 23:50]
      addr <= 64'h0; // @[C2H.scala 23:50]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[C2H.scala 53:39]
        addr <= io_start_addr; // @[C2H.scala 56:65]
      end
    end
    if (reset) begin // @[C2H.scala 24:50]
      length <= 32'h0; // @[C2H.scala 24:50]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[C2H.scala 53:39]
        length <= io_length; // @[C2H.scala 57:65]
      end
    end
    if (reset) begin // @[C2H.scala 25:42]
      valid_cmd <= 1'h0; // @[C2H.scala 25:42]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[C2H.scala 66:48]
          valid_cmd <= 1'h0; // @[C2H.scala 68:65]
        end else begin
          valid_cmd <= 1'h1; // @[C2H.scala 65:65]
        end
      end
    end
    if (reset) begin // @[C2H.scala 29:42]
      count_time <= 32'h0; // @[C2H.scala 29:42]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[C2H.scala 53:39]
        count_time <= 32'h0; // @[C2H.scala 59:65]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      count_time <= _count_time_T_1; // @[C2H.scala 64:65]
    end
    if (reset) begin // @[C2H.scala 30:42]
      send_cmd_count <= 32'h0; // @[C2H.scala 30:42]
    end else if (_T_2) begin // @[C2H.scala 81:32]
      send_cmd_count <= _send_cmd_count_T_1; // @[C2H.scala 82:33]
    end
    complete <= reset | _GEN_21; // @[C2H.scala 33:42 C2H.scala 33:42]
    if (reset) begin // @[C2H.scala 35:50]
      hold <= 4'h0; // @[C2H.scala 35:50]
    end else if (!(_T)) begin // @[Conditional.scala 40:58]
      if (_T_1) begin // @[Conditional.scala 39:67]
        if (_T_2) begin // @[C2H.scala 66:48]
          hold <= 4'ha; // @[C2H.scala 69:65]
        end
      end else if (_T_3) begin // @[Conditional.scala 39:67]
        hold <= _hold_T_1; // @[C2H.scala 73:30]
      end
    end
    if (reset) begin // @[C2H.scala 48:42]
      state_cmd <= 2'h0; // @[C2H.scala 48:42]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[C2H.scala 53:39]
        state_cmd <= 2'h1; // @[C2H.scala 54:65]
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      if (_T_2) begin // @[C2H.scala 66:48]
        state_cmd <= 2'h2; // @[C2H.scala 67:65]
      end
    end else if (_T_3) begin // @[Conditional.scala 39:67]
      state_cmd <= _GEN_11;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addr = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  length = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  valid_cmd = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  count_time = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  send_cmd_count = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  complete = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  hold = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  state_cmd = _RAND_7[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module C2H_Complete(
  input         clock,
  input         reset,
  input  [63:0] io_h2c_cpt_addr,
  input  [63:0] io_c2h_cpt_addr,
  input  [63:0] io_p2p_cpt_addr,
  input         io_h2c_complete,
  input         io_c2h_complete,
  input         io_p2p_complete,
  input  [31:0] io_pfch_tag,
  input         io_h2c_start,
  input         io_c2h_start,
  output        io_h2c_cpt_complete,
  output        io_c2h_cpt_complete,
  output        io_p2p_cpt_complete,
  input  [31:0] io_polling,
  input         io_c2h_cmd_ready,
  output        io_c2h_cmd_valid,
  output [63:0] io_c2h_cmd_bits_addr,
  output [6:0]  io_c2h_cmd_bits_pfch_tag,
  input         io_c2h_data_ready,
  output        io_c2h_data_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  _h2c_cpt_start_T = io_polling == 32'h1; // @[C2H_Complete.scala 33:36]
  reg  h2c_cpt_start_REG; // @[C2H_Complete.scala 33:80]
  wire  h2c_cpt_start = io_polling == 32'h1 & io_h2c_complete & ~h2c_cpt_start_REG; // @[C2H_Complete.scala 33:70]
  reg  c2h_cpt_start_REG; // @[C2H_Complete.scala 34:80]
  wire  c2h_cpt_start = _h2c_cpt_start_T & io_c2h_complete & ~c2h_cpt_start_REG; // @[C2H_Complete.scala 34:70]
  wire  p2p_cpt_start = _h2c_cpt_start_T & io_p2p_complete; // @[C2H_Complete.scala 35:44]
  reg  cmd_valid; // @[C2H_Complete.scala 36:28]
  reg  data_valid; // @[C2H_Complete.scala 37:29]
  reg [63:0] cpt_addr; // @[C2H_Complete.scala 38:27]
  reg [63:0] h2c_cpt_addr; // @[C2H_Complete.scala 39:31]
  reg [63:0] c2h_cpt_addr; // @[C2H_Complete.scala 40:31]
  reg  h2c_cpt_complete; // @[C2H_Complete.scala 42:35]
  reg  c2h_cpt_complete; // @[C2H_Complete.scala 43:35]
  reg  p2p_cpt_complete; // @[C2H_Complete.scala 44:35]
  wire  _GEN_1 = io_h2c_start ? 1'h0 : h2c_cpt_complete; // @[C2H_Complete.scala 50:9 C2H_Complete.scala 52:30 C2H_Complete.scala 42:35]
  wire  _GEN_3 = io_c2h_start ? 1'h0 : c2h_cpt_complete; // @[C2H_Complete.scala 55:9 C2H_Complete.scala 57:30 C2H_Complete.scala 43:35]
  wire  _GEN_4 = p2p_cpt_complete ? 1'h0 : p2p_cpt_complete; // @[C2H_Complete.scala 60:5 C2H_Complete.scala 61:26 C2H_Complete.scala 44:35]
  reg  cmd_fire; // @[C2H_Complete.scala 84:27]
  reg  data_fire; // @[C2H_Complete.scala 85:28]
  reg  p2p_started; // @[C2H_Complete.scala 86:30]
  reg  h2c_started; // @[C2H_Complete.scala 87:30]
  reg  c2h_started; // @[C2H_Complete.scala 88:30]
  wire  _GEN_5 = p2p_cpt_start | cmd_valid; // @[C2H_Complete.scala 92:9 C2H_Complete.scala 93:23 C2H_Complete.scala 36:28]
  wire  _GEN_6 = p2p_cpt_start | data_valid; // @[C2H_Complete.scala 92:9 C2H_Complete.scala 94:24 C2H_Complete.scala 37:29]
  wire  _GEN_8 = p2p_cpt_start | p2p_started; // @[C2H_Complete.scala 92:9 C2H_Complete.scala 96:25 C2H_Complete.scala 86:30]
  wire  _GEN_9 = h2c_cpt_start | _GEN_5; // @[C2H_Complete.scala 100:9 C2H_Complete.scala 101:23]
  wire  _GEN_10 = h2c_cpt_start | _GEN_6; // @[C2H_Complete.scala 100:9 C2H_Complete.scala 102:24]
  wire  _GEN_12 = h2c_cpt_start | h2c_started; // @[C2H_Complete.scala 100:9 C2H_Complete.scala 104:25 C2H_Complete.scala 87:30]
  wire  _GEN_13 = c2h_cpt_start | _GEN_9; // @[C2H_Complete.scala 109:9 C2H_Complete.scala 110:23]
  wire  _GEN_14 = c2h_cpt_start | _GEN_10; // @[C2H_Complete.scala 109:9 C2H_Complete.scala 111:24]
  wire  _GEN_16 = c2h_cpt_start | c2h_started; // @[C2H_Complete.scala 109:9 C2H_Complete.scala 113:25 C2H_Complete.scala 88:30]
  wire  _T = io_c2h_cmd_ready & io_c2h_cmd_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_18 = _T | cmd_fire; // @[C2H_Complete.scala 118:9 C2H_Complete.scala 120:22 C2H_Complete.scala 84:27]
  wire  _T_1 = io_c2h_data_ready & io_c2h_data_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_20 = _T_1 | data_fire; // @[C2H_Complete.scala 123:9 C2H_Complete.scala 125:23 C2H_Complete.scala 85:28]
  wire  _T_2 = cmd_fire & data_fire; // @[C2H_Complete.scala 127:20]
  wire  _GEN_22 = p2p_started | _GEN_4; // @[C2H_Complete.scala 132:13 C2H_Complete.scala 134:34]
  wire  _GEN_24 = h2c_started | _GEN_1; // @[C2H_Complete.scala 137:13 C2H_Complete.scala 139:34]
  wire  _GEN_26 = c2h_started | _GEN_3; // @[C2H_Complete.scala 142:13 C2H_Complete.scala 144:34]
  wire  _GEN_30 = _T_2 ? _GEN_22 : _GEN_4; // @[C2H_Complete.scala 128:9]
  wire  _GEN_32 = _T_2 ? _GEN_24 : _GEN_1; // @[C2H_Complete.scala 128:9]
  wire  _GEN_34 = _T_2 ? _GEN_26 : _GEN_3; // @[C2H_Complete.scala 128:9]
  assign io_h2c_cpt_complete = h2c_cpt_complete; // @[C2H_Complete.scala 45:25]
  assign io_c2h_cpt_complete = c2h_cpt_complete; // @[C2H_Complete.scala 46:25]
  assign io_p2p_cpt_complete = p2p_cpt_complete; // @[C2H_Complete.scala 47:25]
  assign io_c2h_cmd_valid = cmd_valid; // @[C2H_Complete.scala 77:33]
  assign io_c2h_cmd_bits_addr = cpt_addr; // @[C2H_Complete.scala 73:41]
  assign io_c2h_cmd_bits_pfch_tag = io_pfch_tag[6:0]; // @[C2H_Complete.scala 75:33]
  assign io_c2h_data_valid = data_valid; // @[C2H_Complete.scala 80:33]
  always @(posedge clock) begin
    h2c_cpt_start_REG <= io_h2c_complete; // @[C2H_Complete.scala 33:96]
    c2h_cpt_start_REG <= io_c2h_complete; // @[C2H_Complete.scala 34:96]
    if (reset) begin // @[C2H_Complete.scala 36:28]
      cmd_valid <= 1'h0; // @[C2H_Complete.scala 36:28]
    end else if (_T) begin // @[C2H_Complete.scala 118:9]
      cmd_valid <= 1'h0; // @[C2H_Complete.scala 119:23]
    end else begin
      cmd_valid <= _GEN_13;
    end
    if (reset) begin // @[C2H_Complete.scala 37:29]
      data_valid <= 1'h0; // @[C2H_Complete.scala 37:29]
    end else if (_T_1) begin // @[C2H_Complete.scala 123:9]
      data_valid <= 1'h0; // @[C2H_Complete.scala 124:24]
    end else begin
      data_valid <= _GEN_14;
    end
    if (reset) begin // @[C2H_Complete.scala 38:27]
      cpt_addr <= 64'h0; // @[C2H_Complete.scala 38:27]
    end else if (c2h_cpt_start) begin // @[C2H_Complete.scala 109:9]
      cpt_addr <= c2h_cpt_addr; // @[C2H_Complete.scala 112:22]
    end else if (h2c_cpt_start) begin // @[C2H_Complete.scala 100:9]
      cpt_addr <= h2c_cpt_addr; // @[C2H_Complete.scala 103:22]
    end else if (p2p_cpt_start) begin // @[C2H_Complete.scala 92:9]
      cpt_addr <= io_p2p_cpt_addr; // @[C2H_Complete.scala 95:22]
    end
    if (reset) begin // @[C2H_Complete.scala 39:31]
      h2c_cpt_addr <= 64'h0; // @[C2H_Complete.scala 39:31]
    end else if (io_h2c_start) begin // @[C2H_Complete.scala 50:9]
      h2c_cpt_addr <= io_h2c_cpt_addr; // @[C2H_Complete.scala 51:26]
    end
    if (reset) begin // @[C2H_Complete.scala 40:31]
      c2h_cpt_addr <= 64'h0; // @[C2H_Complete.scala 40:31]
    end else if (io_c2h_start) begin // @[C2H_Complete.scala 55:9]
      c2h_cpt_addr <= io_c2h_cpt_addr; // @[C2H_Complete.scala 56:26]
    end
    h2c_cpt_complete <= reset | _GEN_32; // @[C2H_Complete.scala 42:35 C2H_Complete.scala 42:35]
    c2h_cpt_complete <= reset | _GEN_34; // @[C2H_Complete.scala 43:35 C2H_Complete.scala 43:35]
    p2p_cpt_complete <= reset | _GEN_30; // @[C2H_Complete.scala 44:35 C2H_Complete.scala 44:35]
    if (reset) begin // @[C2H_Complete.scala 84:27]
      cmd_fire <= 1'h0; // @[C2H_Complete.scala 84:27]
    end else if (_T_2) begin // @[C2H_Complete.scala 128:9]
      cmd_fire <= 1'h0; // @[C2H_Complete.scala 129:22]
    end else begin
      cmd_fire <= _GEN_18;
    end
    if (reset) begin // @[C2H_Complete.scala 85:28]
      data_fire <= 1'h0; // @[C2H_Complete.scala 85:28]
    end else if (_T_2) begin // @[C2H_Complete.scala 128:9]
      data_fire <= 1'h0; // @[C2H_Complete.scala 130:23]
    end else begin
      data_fire <= _GEN_20;
    end
    if (reset) begin // @[C2H_Complete.scala 86:30]
      p2p_started <= 1'h0; // @[C2H_Complete.scala 86:30]
    end else if (_T_2) begin // @[C2H_Complete.scala 128:9]
      if (p2p_started) begin // @[C2H_Complete.scala 132:13]
        p2p_started <= 1'h0; // @[C2H_Complete.scala 133:29]
      end else begin
        p2p_started <= _GEN_8;
      end
    end else begin
      p2p_started <= _GEN_8;
    end
    if (reset) begin // @[C2H_Complete.scala 87:30]
      h2c_started <= 1'h0; // @[C2H_Complete.scala 87:30]
    end else if (_T_2) begin // @[C2H_Complete.scala 128:9]
      if (h2c_started) begin // @[C2H_Complete.scala 137:13]
        h2c_started <= 1'h0; // @[C2H_Complete.scala 138:29]
      end else begin
        h2c_started <= _GEN_12;
      end
    end else begin
      h2c_started <= _GEN_12;
    end
    if (reset) begin // @[C2H_Complete.scala 88:30]
      c2h_started <= 1'h0; // @[C2H_Complete.scala 88:30]
    end else if (_T_2) begin // @[C2H_Complete.scala 128:9]
      if (c2h_started) begin // @[C2H_Complete.scala 142:13]
        c2h_started <= 1'h0; // @[C2H_Complete.scala 143:29]
      end else begin
        c2h_started <= _GEN_16;
      end
    end else begin
      c2h_started <= _GEN_16;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  h2c_cpt_start_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  c2h_cpt_start_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cmd_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  data_valid = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  cpt_addr = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  h2c_cpt_addr = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  c2h_cpt_addr = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  h2c_cpt_complete = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  c2h_cpt_complete = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  p2p_cpt_complete = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  cmd_fire = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  data_fire = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  p2p_started = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  h2c_started = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  c2h_started = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module H2M(
  input         clock,
  input         reset,
  input  [33:0] io_start_addr,
  input  [31:0] io_length,
  input         io_start,
  output        io_complete,
  output [33:0] io_awaddr,
  output        io_awvalid,
  input         io_awready,
  output [7:0]  io_awlen,
  input         io_wfire,
  output        io_fifo_rden,
  output        io_wlast,
  input         io_last,
  output        io_clear
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[H2M.scala 31:34]
  reg  init; // @[H2M.scala 32:34]
  reg [31:0] length; // @[H2M.scala 34:34]
  reg [31:0] total_length; // @[H2M.scala 35:34]
  reg  complete; // @[H2M.scala 36:34]
  reg [33:0] awaddr; // @[H2M.scala 37:34]
  reg  awvalid; // @[H2M.scala 38:34]
  reg [7:0] awlen; // @[H2M.scala 39:34]
  reg  wlast; // @[H2M.scala 40:34]
  reg  last; // @[H2M.scala 41:34]
  reg  clear; // @[H2M.scala 42:34]
  reg [31:0] write_count; // @[H2M.scala 43:34]
  reg [33:0] end_addr; // @[H2M.scala 45:34]
  reg [33:0] tmp_addr; // @[H2M.scala 46:34]
  reg [33:0] next_addr; // @[H2M.scala 47:34]
  reg [7:0] write_len; // @[H2M.scala 48:34]
  wire [31:0] _write_count_T_1 = write_count + 32'h20; // @[H2M.scala 53:37]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [31:0] _total_length_T_1 = total_length + io_length; // @[H2M.scala 60:49]
  wire [33:0] _GEN_128 = {{2'd0}, io_length}; // @[H2M.scala 64:50]
  wire [33:0] _end_addr_T_1 = io_start_addr + _GEN_128; // @[H2M.scala 64:50]
  wire [31:0] _GEN_129 = {{23'd0}, io_start_addr[8:0]}; // @[H2M.scala 67:50]
  wire [31:0] _T_3 = _GEN_129 + io_length; // @[H2M.scala 67:50]
  wire [24:0] _next_addr_T_2 = io_start_addr[33:9] + 25'h1; // @[H2M.scala 68:59]
  wire [33:0] _next_addr_T_3 = {_next_addr_T_2,9'h0}; // @[Cat.scala 30:58]
  wire [33:0] _GEN_1 = 32'h200 < _T_3 ? _next_addr_T_3 : _end_addr_T_1; // @[H2M.scala 67:62 H2M.scala 68:33 H2M.scala 70:33]
  wire  _GEN_6 = io_start ? 1'h0 : complete; // @[H2M.scala 57:28 H2M.scala 62:33 H2M.scala 36:34]
  wire [24:0] _T_8 = next_addr[33:9] + 25'h1; // @[H2M.scala 82:38]
  wire [33:0] _next_addr_T_7 = next_addr + 34'h200; // @[H2M.scala 83:46]
  wire [33:0] _GEN_14 = _T_8 <= end_addr[33:9] ? _next_addr_T_7 : end_addr; // @[H2M.scala 82:61 H2M.scala 83:33 H2M.scala 85:33]
  wire [33:0] _awlen_T_1 = next_addr - tmp_addr; // @[H2M.scala 88:38]
  wire [3:0] _awlen_T_4 = _awlen_T_1[8:5] - 4'h1; // @[H2M.scala 88:54]
  wire  _GEN_20 = init | awvalid; // @[H2M.scala 73:24 H2M.scala 87:26 H2M.scala 38:34]
  wire  _T_11 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_22 = awvalid & io_awready ? 1'h0 : awvalid; // @[H2M.scala 92:50 H2M.scala 93:29 H2M.scala 38:34]
  wire [1:0] _GEN_23 = awvalid & io_awready ? 2'h2 : state; // @[H2M.scala 92:50 H2M.scala 94:29 H2M.scala 31:34]
  wire [7:0] _write_len_T_1 = write_len + 8'h1; // @[H2M.scala 98:54]
  wire  _T_15 = tmp_addr == end_addr; // @[H2M.scala 100:36]
  wire [1:0] _GEN_25 = tmp_addr == end_addr ? 2'h3 : 2'h1; // @[H2M.scala 100:50 H2M.scala 101:41 H2M.scala 104:41]
  wire [7:0] _GEN_26 = tmp_addr == end_addr ? _write_len_T_1 : 8'h0; // @[H2M.scala 100:50 H2M.scala 98:41 H2M.scala 105:41]
  wire [33:0] _GEN_27 = tmp_addr == end_addr ? awaddr : tmp_addr; // @[H2M.scala 100:50 H2M.scala 37:34 H2M.scala 106:41]
  wire [33:0] _GEN_28 = tmp_addr == end_addr ? tmp_addr : next_addr; // @[H2M.scala 100:50 H2M.scala 46:34 H2M.scala 107:41]
  wire [33:0] _GEN_29 = tmp_addr == end_addr ? next_addr : _GEN_14; // @[H2M.scala 100:50 H2M.scala 47:34]
  wire  _GEN_30 = tmp_addr == end_addr ? _GEN_22 : 1'h1; // @[H2M.scala 100:50 H2M.scala 113:41]
  wire [7:0] _GEN_31 = tmp_addr == end_addr ? awlen : {{4'd0}, _awlen_T_4}; // @[H2M.scala 100:50 H2M.scala 39:34 H2M.scala 114:37]
  wire [1:0] _GEN_32 = awlen == 8'h0 ? _GEN_25 : _GEN_23; // @[H2M.scala 99:38]
  wire [7:0] _GEN_33 = awlen == 8'h0 ? _GEN_26 : _write_len_T_1; // @[H2M.scala 99:38 H2M.scala 98:41]
  wire [33:0] _GEN_34 = awlen == 8'h0 ? _GEN_27 : awaddr; // @[H2M.scala 99:38 H2M.scala 37:34]
  wire [33:0] _GEN_35 = awlen == 8'h0 ? _GEN_28 : tmp_addr; // @[H2M.scala 99:38 H2M.scala 46:34]
  wire [33:0] _GEN_36 = awlen == 8'h0 ? _GEN_29 : next_addr; // @[H2M.scala 99:38 H2M.scala 47:34]
  wire  _GEN_37 = awlen == 8'h0 ? _GEN_30 : _GEN_22; // @[H2M.scala 99:38]
  wire [7:0] _GEN_38 = awlen == 8'h0 ? _GEN_31 : awlen; // @[H2M.scala 99:38 H2M.scala 39:34]
  wire  _T_21 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [7:0] _T_23 = awlen - 8'h1; // @[H2M.scala 121:43]
  wire  _T_24 = write_len == _T_23; // @[H2M.scala 121:33]
  wire  _GEN_53 = _T_15 ? awvalid : 1'h1; // @[H2M.scala 128:50 H2M.scala 38:34 H2M.scala 141:41]
  wire [1:0] _GEN_55 = write_len == awlen ? _GEN_25 : state; // @[H2M.scala 127:44 H2M.scala 31:34]
  wire [7:0] _GEN_56 = write_len == awlen ? _GEN_26 : _write_len_T_1; // @[H2M.scala 127:44 H2M.scala 126:41]
  wire [33:0] _GEN_57 = write_len == awlen ? _GEN_27 : awaddr; // @[H2M.scala 127:44 H2M.scala 37:34]
  wire [33:0] _GEN_58 = write_len == awlen ? _GEN_28 : tmp_addr; // @[H2M.scala 127:44 H2M.scala 46:34]
  wire [33:0] _GEN_59 = write_len == awlen ? _GEN_29 : next_addr; // @[H2M.scala 127:44 H2M.scala 47:34]
  wire  _GEN_60 = write_len == awlen ? _GEN_53 : awvalid; // @[H2M.scala 127:44 H2M.scala 38:34]
  wire [7:0] _GEN_61 = write_len == awlen ? _GEN_31 : awlen; // @[H2M.scala 127:44 H2M.scala 39:34]
  wire  _GEN_62 = io_wfire ? _T_24 : wlast; // @[H2M.scala 120:28 H2M.scala 40:34]
  wire [7:0] _GEN_63 = io_wfire ? _GEN_56 : write_len; // @[H2M.scala 120:28 H2M.scala 48:34]
  wire [1:0] _GEN_64 = io_wfire ? _GEN_55 : state; // @[H2M.scala 120:28 H2M.scala 31:34]
  wire [33:0] _GEN_65 = io_wfire ? _GEN_57 : awaddr; // @[H2M.scala 120:28 H2M.scala 37:34]
  wire [33:0] _GEN_66 = io_wfire ? _GEN_58 : tmp_addr; // @[H2M.scala 120:28 H2M.scala 46:34]
  wire [33:0] _GEN_67 = io_wfire ? _GEN_59 : next_addr; // @[H2M.scala 120:28 H2M.scala 47:34]
  wire  _GEN_68 = io_wfire ? _GEN_60 : awvalid; // @[H2M.scala 120:28 H2M.scala 38:34]
  wire [7:0] _GEN_69 = io_wfire ? _GEN_61 : awlen; // @[H2M.scala 120:28 H2M.scala 39:34]
  wire  _T_32 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_33 = write_count == total_length; // @[H2M.scala 149:35]
  wire [1:0] _GEN_70 = _T_33 ? 2'h0 : state; // @[H2M.scala 150:21 H2M.scala 151:41 H2M.scala 31:34]
  wire [33:0] _GEN_71 = _T_33 ? 34'h0 : awaddr; // @[H2M.scala 150:21 H2M.scala 152:41 H2M.scala 37:34]
  wire  _GEN_72 = _T_33 ? 1'h0 : awvalid; // @[H2M.scala 150:21 H2M.scala 153:41 H2M.scala 38:34]
  wire [7:0] _GEN_73 = _T_33 ? 8'h0 : awlen; // @[H2M.scala 150:21 H2M.scala 154:41 H2M.scala 39:34]
  wire  _GEN_74 = _T_33 ? 1'h0 : wlast; // @[H2M.scala 150:21 H2M.scala 155:41 H2M.scala 40:34]
  wire [7:0] _GEN_75 = _T_33 ? 8'h0 : write_len; // @[H2M.scala 150:21 H2M.scala 157:41 H2M.scala 48:34]
  wire  _GEN_77 = _T_33 | clear; // @[H2M.scala 150:21 H2M.scala 159:41 H2M.scala 42:34]
  wire [1:0] _GEN_78 = last ? _GEN_70 : 2'h0; // @[H2M.scala 148:24 H2M.scala 164:33]
  wire [33:0] _GEN_79 = last ? _GEN_71 : 34'h0; // @[H2M.scala 148:24 H2M.scala 165:33]
  wire  _GEN_80 = last & _GEN_72; // @[H2M.scala 148:24 H2M.scala 166:33]
  wire [7:0] _GEN_81 = last ? _GEN_73 : 8'h0; // @[H2M.scala 148:24 H2M.scala 167:33]
  wire  _GEN_82 = last & _GEN_74; // @[H2M.scala 148:24 H2M.scala 168:33]
  wire [7:0] _GEN_83 = last ? _GEN_75 : 8'h0; // @[H2M.scala 148:24 H2M.scala 170:33]
  wire  _GEN_84 = last ? _T_33 : 1'h1; // @[H2M.scala 148:24 H2M.scala 171:33]
  wire  _GEN_85 = last ? _GEN_77 : clear; // @[H2M.scala 148:24 H2M.scala 42:34]
  wire [1:0] _GEN_86 = _T_32 ? _GEN_78 : state; // @[Conditional.scala 39:67 H2M.scala 31:34]
  wire [33:0] _GEN_87 = _T_32 ? _GEN_79 : awaddr; // @[Conditional.scala 39:67 H2M.scala 37:34]
  wire  _GEN_88 = _T_32 ? _GEN_80 : awvalid; // @[Conditional.scala 39:67 H2M.scala 38:34]
  wire [7:0] _GEN_89 = _T_32 ? _GEN_81 : awlen; // @[Conditional.scala 39:67 H2M.scala 39:34]
  wire  _GEN_90 = _T_32 ? _GEN_82 : wlast; // @[Conditional.scala 39:67 H2M.scala 40:34]
  wire [7:0] _GEN_91 = _T_32 ? _GEN_83 : write_len; // @[Conditional.scala 39:67 H2M.scala 48:34]
  wire  _GEN_92 = _T_32 ? _GEN_84 : complete; // @[Conditional.scala 39:67 H2M.scala 36:34]
  wire  _GEN_93 = _T_32 ? _GEN_85 : clear; // @[Conditional.scala 39:67 H2M.scala 42:34]
  wire  _GEN_102 = _T_21 ? complete : _GEN_92; // @[Conditional.scala 39:67 H2M.scala 36:34]
  wire  _GEN_112 = _T_11 ? complete : _GEN_102; // @[Conditional.scala 39:67 H2M.scala 36:34]
  wire  _GEN_118 = _T ? _GEN_6 : _GEN_112; // @[Conditional.scala 40:58]
  wire [10:0] _io_awlen_T = {3'h0,awlen}; // @[Cat.scala 30:58]
  assign io_complete = complete; // @[H2M.scala 180:29]
  assign io_awaddr = awaddr; // @[H2M.scala 176:29]
  assign io_awvalid = awvalid; // @[H2M.scala 177:29]
  assign io_awlen = _io_awlen_T[7:0]; // @[H2M.scala 178:29]
  assign io_fifo_rden = state == 2'h2; // @[H2M.scala 50:35]
  assign io_wlast = wlast; // @[H2M.scala 179:29]
  assign io_clear = clear; // @[H2M.scala 181:29]
  always @(posedge clock) begin
    if (reset) begin // @[H2M.scala 31:34]
      state <= 2'h0; // @[H2M.scala 31:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[H2M.scala 73:24]
        if (length == 32'h0) begin // @[H2M.scala 74:39]
          state <= 2'h3; // @[H2M.scala 75:33]
        end else begin
          state <= 2'h1; // @[H2M.scala 77:33]
        end
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (io_wfire) begin // @[H2M.scala 97:28]
        state <= _GEN_32;
      end else begin
        state <= _GEN_23;
      end
    end else if (_T_21) begin // @[Conditional.scala 39:67]
      state <= _GEN_64;
    end else begin
      state <= _GEN_86;
    end
    init <= io_start; // @[H2M.scala 32:34]
    if (reset) begin // @[H2M.scala 34:34]
      length <= 32'h0; // @[H2M.scala 34:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2M.scala 57:28]
        length <= io_length; // @[H2M.scala 61:33]
      end
    end
    if (reset) begin // @[H2M.scala 35:34]
      total_length <= 32'h0; // @[H2M.scala 35:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2M.scala 57:28]
        total_length <= _total_length_T_1; // @[H2M.scala 60:33]
      end
    end
    complete <= reset | _GEN_118; // @[H2M.scala 36:34 H2M.scala 36:34]
    if (reset) begin // @[H2M.scala 37:34]
      awaddr <= 34'h0; // @[H2M.scala 37:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[H2M.scala 73:24]
        awaddr <= tmp_addr; // @[H2M.scala 80:33]
      end else if (io_start) begin // @[H2M.scala 57:28]
        awaddr <= io_start_addr; // @[H2M.scala 66:33]
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (io_wfire) begin // @[H2M.scala 97:28]
        awaddr <= _GEN_34;
      end
    end else if (_T_21) begin // @[Conditional.scala 39:67]
      awaddr <= _GEN_65;
    end else begin
      awaddr <= _GEN_87;
    end
    if (reset) begin // @[H2M.scala 38:34]
      awvalid <= 1'h0; // @[H2M.scala 38:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      awvalid <= _GEN_20;
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (io_wfire) begin // @[H2M.scala 97:28]
        awvalid <= _GEN_37;
      end else begin
        awvalid <= _GEN_22;
      end
    end else if (_T_21) begin // @[Conditional.scala 39:67]
      awvalid <= _GEN_68;
    end else begin
      awvalid <= _GEN_88;
    end
    if (reset) begin // @[H2M.scala 39:34]
      awlen <= 8'h0; // @[H2M.scala 39:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[H2M.scala 73:24]
        awlen <= {{4'd0}, _awlen_T_4}; // @[H2M.scala 88:25]
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (io_wfire) begin // @[H2M.scala 97:28]
        awlen <= _GEN_38;
      end
    end else if (_T_21) begin // @[Conditional.scala 39:67]
      awlen <= _GEN_69;
    end else begin
      awlen <= _GEN_89;
    end
    if (reset) begin // @[H2M.scala 40:34]
      wlast <= 1'h0; // @[H2M.scala 40:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2M.scala 57:28]
        wlast <= 1'h0; // @[H2M.scala 63:33]
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (_T_21) begin // @[Conditional.scala 39:67]
        wlast <= _GEN_62;
      end else begin
        wlast <= _GEN_90;
      end
    end
    if (reset) begin // @[H2M.scala 41:34]
      last <= 1'h0; // @[H2M.scala 41:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2M.scala 57:28]
        last <= io_last; // @[H2M.scala 59:33]
      end
    end
    if (reset) begin // @[H2M.scala 42:34]
      clear <= 1'h0; // @[H2M.scala 42:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2M.scala 57:28]
        clear <= 1'h0; // @[H2M.scala 58:33]
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (!(_T_21)) begin // @[Conditional.scala 39:67]
        clear <= _GEN_93;
      end
    end
    if (reset) begin // @[H2M.scala 43:34]
      write_count <= 32'h0; // @[H2M.scala 43:34]
    end else if (io_wfire) begin // @[H2M.scala 53:9]
      write_count <= _write_count_T_1; // @[H2M.scala 53:22]
    end
    if (reset) begin // @[H2M.scala 45:34]
      end_addr <= 34'h0; // @[H2M.scala 45:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[H2M.scala 57:28]
        end_addr <= _end_addr_T_1; // @[H2M.scala 64:33]
      end
    end
    if (reset) begin // @[H2M.scala 46:34]
      tmp_addr <= 34'h0; // @[H2M.scala 46:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[H2M.scala 73:24]
        tmp_addr <= next_addr; // @[H2M.scala 81:33]
      end else if (io_start) begin // @[H2M.scala 57:28]
        tmp_addr <= io_start_addr; // @[H2M.scala 65:33]
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (io_wfire) begin // @[H2M.scala 97:28]
        tmp_addr <= _GEN_35;
      end
    end else if (_T_21) begin // @[Conditional.scala 39:67]
      tmp_addr <= _GEN_66;
    end
    if (reset) begin // @[H2M.scala 47:34]
      next_addr <= 34'h0; // @[H2M.scala 47:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[H2M.scala 73:24]
        if (_T_8 <= end_addr[33:9]) begin // @[H2M.scala 82:61]
          next_addr <= _next_addr_T_7; // @[H2M.scala 83:33]
        end else begin
          next_addr <= end_addr; // @[H2M.scala 85:33]
        end
      end else if (io_start) begin // @[H2M.scala 57:28]
        next_addr <= _GEN_1;
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (io_wfire) begin // @[H2M.scala 97:28]
        next_addr <= _GEN_36;
      end
    end else if (_T_21) begin // @[Conditional.scala 39:67]
      next_addr <= _GEN_67;
    end
    if (reset) begin // @[H2M.scala 48:34]
      write_len <= 8'h0; // @[H2M.scala 48:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[H2M.scala 73:24]
        if (!(length == 32'h0)) begin // @[H2M.scala 74:39]
          write_len <= 8'h0; // @[H2M.scala 78:33]
        end
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (io_wfire) begin // @[H2M.scala 97:28]
        write_len <= _GEN_33;
      end
    end else if (_T_21) begin // @[Conditional.scala 39:67]
      write_len <= _GEN_63;
    end else begin
      write_len <= _GEN_91;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  init = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  length = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  total_length = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  complete = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  awaddr = _RAND_5[33:0];
  _RAND_6 = {1{`RANDOM}};
  awvalid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  awlen = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  wlast = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  last = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  clear = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  write_count = _RAND_11[31:0];
  _RAND_12 = {2{`RANDOM}};
  end_addr = _RAND_12[33:0];
  _RAND_13 = {2{`RANDOM}};
  tmp_addr = _RAND_13[33:0];
  _RAND_14 = {2{`RANDOM}};
  next_addr = _RAND_14[33:0];
  _RAND_15 = {1{`RANDOM}};
  write_len = _RAND_15[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module M2H(
  input         clock,
  input         reset,
  input  [33:0] io_start_addr,
  input  [31:0] io_length,
  input         io_start,
  output        io_complete,
  output [33:0] io_araddr,
  output        io_arvalid,
  input         io_arready,
  output [7:0]  io_arlen,
  input         io_rfire,
  input         io_last,
  input         io_m2h_queue_empty,
  input         io_m2h_valid_tmpreg,
  output        io_read_count_equal
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[M2H.scala 31:34]
  reg  init; // @[M2H.scala 32:34]
  reg [31:0] length; // @[M2H.scala 34:34]
  reg [31:0] total_length; // @[M2H.scala 35:34]
  reg  complete; // @[M2H.scala 36:34]
  reg [33:0] araddr; // @[M2H.scala 37:34]
  reg  arvalid; // @[M2H.scala 38:34]
  reg [7:0] arlen; // @[M2H.scala 39:34]
  reg [31:0] read_count; // @[M2H.scala 40:34]
  reg [3:0] hold1; // @[M2H.scala 41:34]
  reg [3:0] hold2; // @[M2H.scala 42:34]
  reg [33:0] end_addr; // @[M2H.scala 44:34]
  reg [33:0] tmp_addr; // @[M2H.scala 45:34]
  reg [33:0] next_addr; // @[M2H.scala 46:34]
  wire [31:0] _read_count_T_1 = read_count + 32'h20; // @[M2H.scala 51:35]
  wire  _io_read_count_equal_T = read_count == total_length; // @[M2H.scala 52:40]
  wire  _T = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [31:0] _total_length_T_1 = total_length + io_length; // @[M2H.scala 57:49]
  wire [33:0] _GEN_72 = {{2'd0}, io_length}; // @[M2H.scala 63:50]
  wire [33:0] _end_addr_T_1 = io_start_addr + _GEN_72; // @[M2H.scala 63:50]
  wire [31:0] _GEN_73 = {{23'd0}, io_start_addr[8:0]}; // @[M2H.scala 66:50]
  wire [31:0] _T_3 = _GEN_73 + io_length; // @[M2H.scala 66:50]
  wire [24:0] _next_addr_T_2 = io_start_addr[33:9] + 25'h1; // @[M2H.scala 67:59]
  wire [33:0] _next_addr_T_3 = {_next_addr_T_2,9'h0}; // @[Cat.scala 30:58]
  wire [33:0] _GEN_1 = 32'h200 < _T_3 ? _next_addr_T_3 : _end_addr_T_1; // @[M2H.scala 66:62 M2H.scala 67:33 M2H.scala 69:33]
  wire  _GEN_7 = io_start ? 1'h0 : complete; // @[M2H.scala 56:28 M2H.scala 62:33 M2H.scala 36:34]
  wire [24:0] _T_7 = next_addr[33:9] + 25'h1; // @[M2H.scala 78:38]
  wire [33:0] _next_addr_T_7 = next_addr + 34'h200; // @[M2H.scala 79:46]
  wire [33:0] _GEN_11 = _T_7 <= end_addr[33:9] ? _next_addr_T_7 : end_addr; // @[M2H.scala 78:61 M2H.scala 79:33 M2H.scala 81:33]
  wire [33:0] _arlen_T_1 = next_addr - tmp_addr; // @[M2H.scala 83:42]
  wire [3:0] _arlen_T_4 = _arlen_T_1[8:5] - 4'h1; // @[M2H.scala 83:58]
  wire  _GEN_18 = init | arvalid; // @[M2H.scala 74:13 M2H.scala 85:33 M2H.scala 38:34]
  wire  _T_11 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_20 = tmp_addr == end_addr ? 1'h0 : arvalid; // @[M2H.scala 99:46 M2H.scala 100:33 M2H.scala 38:34]
  wire [1:0] _GEN_21 = tmp_addr == end_addr ? 2'h3 : state; // @[M2H.scala 99:46 M2H.scala 101:33 M2H.scala 31:34]
  wire  _T_20 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_23 = _io_read_count_equal_T & hold1 != 4'h0; // @[M2H.scala 107:51]
  wire [3:0] _hold1_T_1 = hold1 - 4'h1; // @[M2H.scala 109:40]
  wire [3:0] _GEN_28 = _T_23 ? _hold1_T_1 : hold1; // @[M2H.scala 108:21 M2H.scala 109:31 M2H.scala 41:34]
  wire  _T_27 = hold1 == 4'h0 & io_m2h_queue_empty & hold2 != 4'h0; // @[M2H.scala 111:58]
  wire [3:0] _hold2_T_1 = hold2 - 4'h1; // @[M2H.scala 113:40]
  wire [3:0] _GEN_29 = _T_27 ? _hold2_T_1 : hold2; // @[M2H.scala 112:21 M2H.scala 113:31 M2H.scala 42:34]
  wire  _T_30 = hold2 == 4'h0 & ~io_m2h_valid_tmpreg; // @[M2H.scala 115:37]
  wire [1:0] _GEN_31 = _T_30 ? 2'h0 : state; // @[M2H.scala 116:21 M2H.scala 118:37 M2H.scala 31:34]
  wire [33:0] _GEN_32 = _T_30 ? 34'h0 : araddr; // @[M2H.scala 116:21 M2H.scala 119:37 M2H.scala 37:34]
  wire  _GEN_33 = _T_30 ? 1'h0 : arvalid; // @[M2H.scala 116:21 M2H.scala 120:37 M2H.scala 38:34]
  wire [7:0] _GEN_34 = _T_30 ? 8'h0 : arlen; // @[M2H.scala 116:21 M2H.scala 121:37 M2H.scala 39:34]
  wire [3:0] _GEN_35 = io_last ? _GEN_28 : hold1; // @[M2H.scala 106:27 M2H.scala 41:34]
  wire [3:0] _GEN_36 = io_last ? _GEN_29 : hold2; // @[M2H.scala 106:27 M2H.scala 42:34]
  wire  _GEN_37 = io_last ? _T_30 : 1'h1; // @[M2H.scala 106:27 M2H.scala 126:37]
  wire [1:0] _GEN_38 = io_last ? _GEN_31 : 2'h0; // @[M2H.scala 106:27 M2H.scala 127:37]
  wire [33:0] _GEN_39 = io_last ? _GEN_32 : 34'h0; // @[M2H.scala 106:27 M2H.scala 128:37]
  wire  _GEN_40 = io_last & _GEN_33; // @[M2H.scala 106:27 M2H.scala 129:37]
  wire [7:0] _GEN_41 = io_last ? _GEN_34 : 8'h0; // @[M2H.scala 106:27 M2H.scala 130:37]
  wire  _GEN_44 = _T_20 ? _GEN_37 : complete; // @[Conditional.scala 39:67 M2H.scala 36:34]
  wire  _GEN_57 = _T_11 ? complete : _GEN_44; // @[Conditional.scala 39:67 M2H.scala 36:34]
  wire  _GEN_63 = _T ? _GEN_7 : _GEN_57; // @[Conditional.scala 40:58]
  wire [10:0] _io_arlen_T = {3'h0,arlen}; // @[Cat.scala 30:58]
  assign io_complete = complete; // @[M2H.scala 139:29]
  assign io_araddr = araddr; // @[M2H.scala 136:29]
  assign io_arvalid = arvalid; // @[M2H.scala 137:29]
  assign io_arlen = _io_arlen_T[7:0]; // @[M2H.scala 138:29]
  assign io_read_count_equal = read_count == total_length; // @[M2H.scala 52:40]
  always @(posedge clock) begin
    if (reset) begin // @[M2H.scala 31:34]
      state <= 2'h0; // @[M2H.scala 31:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[M2H.scala 74:13]
        if (length == 32'h0) begin // @[M2H.scala 84:39]
          state <= 2'h3; // @[M2H.scala 84:46]
        end else begin
          state <= 2'h1; // @[M2H.scala 84:76]
        end
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (arvalid & io_arready) begin // @[M2H.scala 89:50]
        state <= _GEN_21;
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67]
      state <= _GEN_38;
    end
    init <= io_start; // @[M2H.scala 32:34]
    if (reset) begin // @[M2H.scala 34:34]
      length <= 32'h0; // @[M2H.scala 34:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[M2H.scala 56:28]
        length <= io_length; // @[M2H.scala 58:33]
      end
    end
    if (reset) begin // @[M2H.scala 35:34]
      total_length <= 32'h0; // @[M2H.scala 35:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[M2H.scala 56:28]
        total_length <= _total_length_T_1; // @[M2H.scala 57:33]
      end
    end
    complete <= reset | _GEN_63; // @[M2H.scala 36:34 M2H.scala 36:34]
    if (reset) begin // @[M2H.scala 37:34]
      araddr <= 34'h0; // @[M2H.scala 37:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[M2H.scala 74:13]
        araddr <= tmp_addr; // @[M2H.scala 76:33]
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (arvalid & io_arready) begin // @[M2H.scala 89:50]
        araddr <= tmp_addr; // @[M2H.scala 91:33]
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67]
      araddr <= _GEN_39;
    end
    if (reset) begin // @[M2H.scala 38:34]
      arvalid <= 1'h0; // @[M2H.scala 38:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      arvalid <= _GEN_18;
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (arvalid & io_arready) begin // @[M2H.scala 89:50]
        arvalid <= _GEN_20;
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67]
      arvalid <= _GEN_40;
    end
    if (reset) begin // @[M2H.scala 39:34]
      arlen <= 8'h0; // @[M2H.scala 39:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[M2H.scala 74:13]
        arlen <= {{4'd0}, _arlen_T_4}; // @[M2H.scala 83:29]
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (arvalid & io_arready) begin // @[M2H.scala 89:50]
        arlen <= {{4'd0}, _arlen_T_4}; // @[M2H.scala 98:29]
      end
    end else if (_T_20) begin // @[Conditional.scala 39:67]
      arlen <= _GEN_41;
    end
    if (reset) begin // @[M2H.scala 40:34]
      read_count <= 32'h0; // @[M2H.scala 40:34]
    end else if (io_rfire) begin // @[M2H.scala 51:9]
      read_count <= _read_count_T_1; // @[M2H.scala 51:21]
    end
    if (reset) begin // @[M2H.scala 41:34]
      hold1 <= 4'ha; // @[M2H.scala 41:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[M2H.scala 56:28]
        hold1 <= 4'ha; // @[M2H.scala 60:33]
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (_T_20) begin // @[Conditional.scala 39:67]
        hold1 <= _GEN_35;
      end
    end
    if (reset) begin // @[M2H.scala 42:34]
      hold2 <= 4'h5; // @[M2H.scala 42:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[M2H.scala 56:28]
        hold2 <= 4'h5; // @[M2H.scala 61:33]
      end
    end else if (!(_T_11)) begin // @[Conditional.scala 39:67]
      if (_T_20) begin // @[Conditional.scala 39:67]
        hold2 <= _GEN_36;
      end
    end
    if (reset) begin // @[M2H.scala 44:34]
      end_addr <= 34'h0; // @[M2H.scala 44:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (io_start) begin // @[M2H.scala 56:28]
        end_addr <= _end_addr_T_1; // @[M2H.scala 63:33]
      end
    end
    if (reset) begin // @[M2H.scala 45:34]
      tmp_addr <= 34'h0; // @[M2H.scala 45:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[M2H.scala 74:13]
        tmp_addr <= next_addr; // @[M2H.scala 75:33]
      end else if (io_start) begin // @[M2H.scala 56:28]
        tmp_addr <= io_start_addr; // @[M2H.scala 64:33]
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (arvalid & io_arready) begin // @[M2H.scala 89:50]
        tmp_addr <= next_addr; // @[M2H.scala 90:33]
      end
    end
    if (reset) begin // @[M2H.scala 46:34]
      next_addr <= 34'h0; // @[M2H.scala 46:34]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (init) begin // @[M2H.scala 74:13]
        next_addr <= _GEN_11;
      end else if (io_start) begin // @[M2H.scala 56:28]
        next_addr <= _GEN_1;
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (arvalid & io_arready) begin // @[M2H.scala 89:50]
        next_addr <= _GEN_11;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  init = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  length = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  total_length = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  complete = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  araddr = _RAND_5[33:0];
  _RAND_6 = {1{`RANDOM}};
  arvalid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  arlen = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  read_count = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  hold1 = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  hold2 = _RAND_10[3:0];
  _RAND_11 = {2{`RANDOM}};
  end_addr = _RAND_11[33:0];
  _RAND_12 = {2{`RANDOM}};
  tmp_addr = _RAND_12[33:0];
  _RAND_13 = {2{`RANDOM}};
  next_addr = _RAND_13[33:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_4(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [66:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [66:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [95:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [66:0] ram [0:15]; // @[Decoupled.scala 218:16]
  wire [66:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 218:16]
  wire [66:0] ram_MPORT_data; // @[Decoupled.scala 218:16]
  wire [3:0] ram_MPORT_addr; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_mask; // @[Decoupled.scala 218:16]
  wire  ram_MPORT_en; // @[Decoupled.scala 218:16]
  reg [3:0] enq_ptr_value; // @[Counter.scala 60:40]
  reg [3:0] deq_ptr_value; // @[Counter.scala 60:40]
  reg  maybe_full; // @[Decoupled.scala 221:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 223:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 224:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 225:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _value_T_1 = enq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  wire [3:0] _value_T_3 = deq_ptr_value + 4'h1; // @[Counter.scala 76:24]
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 218:16]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 241:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 240:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 242:15]
  always @(posedge clock) begin
    if(ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 218:16]
    end
    if (reset) begin // @[Counter.scala 60:40]
      enq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_enq) begin // @[Decoupled.scala 229:17]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Counter.scala 60:40]
      deq_ptr_value <= 4'h0; // @[Counter.scala 60:40]
    end else if (do_deq) begin // @[Decoupled.scala 233:17]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 76:15]
    end
    if (reset) begin // @[Decoupled.scala 221:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 221:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 236:28]
      maybe_full <= do_enq; // @[Decoupled.scala 237:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {3{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[66:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module XQueue_34(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [66:0] io_in_bits,
  input         io_out_ready,
  output        io_out_valid,
  output [66:0] io_out_bits
);
  wire  q_clock; // @[XQueue.scala 85:39]
  wire  q_reset; // @[XQueue.scala 85:39]
  wire  q_io_enq_ready; // @[XQueue.scala 85:39]
  wire  q_io_enq_valid; // @[XQueue.scala 85:39]
  wire [66:0] q_io_enq_bits; // @[XQueue.scala 85:39]
  wire  q_io_deq_ready; // @[XQueue.scala 85:39]
  wire  q_io_deq_valid; // @[XQueue.scala 85:39]
  wire [66:0] q_io_deq_bits; // @[XQueue.scala 85:39]
  Queue_4 q ( // @[XQueue.scala 85:39]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits(q_io_enq_bits),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits(q_io_deq_bits)
  );
  assign io_in_ready = q_io_enq_ready; // @[XQueue.scala 87:34]
  assign io_out_valid = q_io_deq_valid; // @[XQueue.scala 88:34]
  assign io_out_bits = q_io_deq_bits; // @[XQueue.scala 88:34]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = io_in_valid; // @[XQueue.scala 87:34]
  assign q_io_enq_bits = io_in_bits; // @[XQueue.scala 87:34]
  assign q_io_deq_ready = io_out_ready; // @[XQueue.scala 88:34]
endmodule
module h2mcmdbufferready(
  input   clock,
  input   reset,
  output  io_ready,
  input   io_valid,
  input   io_complete
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  ready; // @[h2mcmdbufferready.scala 14:24]
  reg  hold; // @[h2mcmdbufferready.scala 15:24]
  wire  _GEN_0 = hold & io_complete; // @[h2mcmdbufferready.scala 19:5 h2mcmdbufferready.scala 20:15 h2mcmdbufferready.scala 22:15]
  wire  _T = io_ready & io_valid; // @[h2mcmdbufferready.scala 25:20]
  wire  _GEN_2 = _T ? 1'h0 : hold; // @[h2mcmdbufferready.scala 26:5 h2mcmdbufferready.scala 28:14 h2mcmdbufferready.scala 15:24]
  reg  REG; // @[h2mcmdbufferready.scala 31:34]
  wire  _T_2 = io_complete & ~REG; // @[h2mcmdbufferready.scala 31:23]
  wire  _GEN_3 = _T_2 | _GEN_2; // @[h2mcmdbufferready.scala 32:5 h2mcmdbufferready.scala 33:14]
  assign io_ready = ready; // @[h2mcmdbufferready.scala 16:14]
  always @(posedge clock) begin
    if (reset) begin // @[h2mcmdbufferready.scala 14:24]
      ready <= 1'h0; // @[h2mcmdbufferready.scala 14:24]
    end else if (_T) begin // @[h2mcmdbufferready.scala 26:5]
      ready <= 1'h0; // @[h2mcmdbufferready.scala 27:15]
    end else begin
      ready <= _GEN_0;
    end
    hold <= reset | _GEN_3; // @[h2mcmdbufferready.scala 15:24 h2mcmdbufferready.scala 15:24]
    REG <= io_complete; // @[h2mcmdbufferready.scala 31:34]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ready = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hold = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  REG = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module c2h_status(
  input         clock,
  input         reset,
  input         io_c2h_start,
  input         io_c2h_status_last,
  input         io_c2h_status_cmp,
  input         io_c2h_status_valid,
  input         io_c2h_status_error,
  input         io_c2h_status_drop,
  output [31:0] io_c2h_status_last_count,
  output [31:0] io_c2h_status_cmp_count,
  output [31:0] io_c2h_status_valid_count,
  output [31:0] io_c2h_status_error_count,
  output [31:0] io_c2h_status_drop_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] c2h_status_last_count; // @[c2hstatus.scala 22:42]
  reg [31:0] c2h_status_cmp_count; // @[c2hstatus.scala 23:42]
  reg [31:0] c2h_status_valid_count; // @[c2hstatus.scala 24:42]
  reg [31:0] c2h_status_error_count; // @[c2hstatus.scala 25:42]
  reg [31:0] c2h_status_drop_count; // @[c2hstatus.scala 26:42]
  wire  _T_3 = io_c2h_status_last & io_c2h_status_valid; // @[c2hstatus.scala 36:38]
  wire [31:0] _c2h_status_last_count_T_1 = c2h_status_last_count + 32'h1; // @[c2hstatus.scala 37:57]
  wire  _T_6 = io_c2h_status_cmp & io_c2h_status_valid; // @[c2hstatus.scala 38:37]
  wire [31:0] _c2h_status_cmp_count_T_1 = c2h_status_cmp_count + 32'h1; // @[c2hstatus.scala 39:55]
  wire [31:0] _c2h_status_valid_count_T_1 = c2h_status_valid_count + 32'h1; // @[c2hstatus.scala 41:59]
  wire  _T_10 = io_c2h_status_error & io_c2h_status_valid; // @[c2hstatus.scala 42:39]
  wire [31:0] _c2h_status_error_count_T_1 = c2h_status_error_count + 32'h1; // @[c2hstatus.scala 43:59]
  wire  _T_13 = io_c2h_status_drop & io_c2h_status_valid; // @[c2hstatus.scala 44:38]
  wire [31:0] _c2h_status_drop_count_T_1 = c2h_status_drop_count + 32'h1; // @[c2hstatus.scala 45:57]
  assign io_c2h_status_last_count = c2h_status_last_count; // @[c2hstatus.scala 46:30]
  assign io_c2h_status_cmp_count = c2h_status_cmp_count; // @[c2hstatus.scala 47:29]
  assign io_c2h_status_valid_count = c2h_status_valid_count; // @[c2hstatus.scala 48:31]
  assign io_c2h_status_error_count = c2h_status_error_count; // @[c2hstatus.scala 49:31]
  assign io_c2h_status_drop_count = c2h_status_drop_count; // @[c2hstatus.scala 50:30]
  always @(posedge clock) begin
    if (reset) begin // @[c2hstatus.scala 22:42]
      c2h_status_last_count <= 32'h0; // @[c2hstatus.scala 22:42]
    end else if (_T_3) begin // @[c2hstatus.scala 37:9]
      c2h_status_last_count <= _c2h_status_last_count_T_1; // @[c2hstatus.scala 37:32]
    end else if (io_c2h_start) begin // @[c2hstatus.scala 28:32]
      c2h_status_last_count <= 32'h0; // @[c2hstatus.scala 29:33]
    end
    if (reset) begin // @[c2hstatus.scala 23:42]
      c2h_status_cmp_count <= 32'h0; // @[c2hstatus.scala 23:42]
    end else if (_T_6) begin // @[c2hstatus.scala 39:9]
      c2h_status_cmp_count <= _c2h_status_cmp_count_T_1; // @[c2hstatus.scala 39:31]
    end else if (io_c2h_start) begin // @[c2hstatus.scala 28:32]
      c2h_status_cmp_count <= 32'h0; // @[c2hstatus.scala 30:33]
    end
    if (reset) begin // @[c2hstatus.scala 24:42]
      c2h_status_valid_count <= 32'h0; // @[c2hstatus.scala 24:42]
    end else if (io_c2h_status_valid) begin // @[c2hstatus.scala 41:9]
      c2h_status_valid_count <= _c2h_status_valid_count_T_1; // @[c2hstatus.scala 41:33]
    end else if (io_c2h_start) begin // @[c2hstatus.scala 28:32]
      c2h_status_valid_count <= 32'h0; // @[c2hstatus.scala 31:33]
    end
    if (reset) begin // @[c2hstatus.scala 25:42]
      c2h_status_error_count <= 32'h0; // @[c2hstatus.scala 25:42]
    end else if (_T_10) begin // @[c2hstatus.scala 43:9]
      c2h_status_error_count <= _c2h_status_error_count_T_1; // @[c2hstatus.scala 43:33]
    end else if (io_c2h_start) begin // @[c2hstatus.scala 28:32]
      c2h_status_error_count <= 32'h0; // @[c2hstatus.scala 32:33]
    end
    if (reset) begin // @[c2hstatus.scala 26:42]
      c2h_status_drop_count <= 32'h0; // @[c2hstatus.scala 26:42]
    end else if (_T_13) begin // @[c2hstatus.scala 45:9]
      c2h_status_drop_count <= _c2h_status_drop_count_T_1; // @[c2hstatus.scala 45:32]
    end else if (io_c2h_start) begin // @[c2hstatus.scala 28:32]
      c2h_status_drop_count <= 32'h0; // @[c2hstatus.scala 33:33]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c2h_status_last_count = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  c2h_status_cmp_count = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2h_status_valid_count = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  c2h_status_error_count = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  c2h_status_drop_count = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module validreg(
  input   clock,
  input   reset,
  input   io_ready,
  input   io_valid,
  output  io_tmpreg
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  tmpreg; // @[validreg.scala 17:26]
  wire  _T_2 = io_valid & ~io_ready; // @[validreg.scala 20:27]
  wire  _GEN_0 = _T_2 | tmpreg; // @[validreg.scala 21:9 validreg.scala 21:17 validreg.scala 17:26]
  wire  _T_5 = tmpreg & io_ready; // @[validreg.scala 23:25]
  assign io_tmpreg = tmpreg; // @[validreg.scala 26:15]
  always @(posedge clock) begin
    if (reset) begin // @[validreg.scala 17:26]
      tmpreg <= 1'h0; // @[validreg.scala 17:26]
    end else if (_T_5) begin // @[validreg.scala 24:9]
      tmpreg <= 1'h0; // @[validreg.scala 24:17]
    end else begin
      tmpreg <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tmpreg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module p2p_counter(
  input         clock,
  input         reset,
  input         io_start,
  input  [31:0] io_length,
  input         io_wready,
  input         io_wvalid,
  input  [31:0] io_wdatasample,
  output        io_p2p_complete,
  input         io_p2p_cpt_complete
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] counter; // @[p2p_counter.scala 24:27]
  wire  _T_4 = io_start & io_wready & io_wvalid & io_wdatasample == 32'hffffffff; // @[p2p_counter.scala 25:44]
  wire [31:0] _counter_T_1 = counter + 32'h20; // @[p2p_counter.scala 27:28]
  reg [31:0] length; // @[p2p_counter.scala 29:25]
  reg  p2p_complete; // @[p2p_counter.scala 31:31]
  reg  working; // @[p2p_counter.scala 32:26]
  wire  _T_6 = working & counter == length; // @[p2p_counter.scala 47:19]
  wire  _GEN_5 = _T_6 | p2p_complete; // @[p2p_counter.scala 48:5 p2p_counter.scala 49:22 p2p_counter.scala 31:31]
  wire  _T_7 = io_p2p_cpt_complete & p2p_complete; // @[p2p_counter.scala 53:31]
  assign io_p2p_complete = p2p_complete; // @[p2p_counter.scala 33:21]
  always @(posedge clock) begin
    if (reset) begin // @[p2p_counter.scala 24:27]
      counter <= 32'h0; // @[p2p_counter.scala 24:27]
    end else if (_T_6) begin // @[p2p_counter.scala 48:5]
      counter <= 32'h0; // @[p2p_counter.scala 50:21]
    end else if (io_start) begin // @[p2p_counter.scala 37:5]
      if (_T_4) begin // @[p2p_counter.scala 26:5]
        counter <= _counter_T_1; // @[p2p_counter.scala 27:17]
      end
    end else begin
      counter <= 32'h0; // @[p2p_counter.scala 44:21]
    end
    if (reset) begin // @[p2p_counter.scala 29:25]
      length <= 32'h0; // @[p2p_counter.scala 29:25]
    end else if (io_start) begin // @[p2p_counter.scala 37:5]
      length <= io_length; // @[p2p_counter.scala 38:21]
    end
    if (reset) begin // @[p2p_counter.scala 31:31]
      p2p_complete <= 1'h0; // @[p2p_counter.scala 31:31]
    end else if (_T_7) begin // @[p2p_counter.scala 54:5]
      p2p_complete <= 1'h0; // @[p2p_counter.scala 55:22]
    end else begin
      p2p_complete <= _GEN_5;
    end
    if (reset) begin // @[p2p_counter.scala 32:26]
      working <= 1'h0; // @[p2p_counter.scala 32:26]
    end else begin
      working <= io_start;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  length = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  p2p_complete = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  working = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  output [15:0] qdma_pin_tx_p,
  output [15:0] qdma_pin_tx_n,
  input  [15:0] qdma_pin_rx_p,
  input  [15:0] qdma_pin_rx_n,
  input         qdma_pin_sys_clk_p,
  input         qdma_pin_sys_clk_n,
  input         qdma_pin_sys_rst_n,
  input         sys_100M_0_p,
  input         sys_100M_0_n
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire  mmcm_io_CLKIN1; // @[Top.scala 16:26]
  wire  mmcm_io_LOCKED; // @[Top.scala 16:26]
  wire  mmcm_io_CLKOUT0; // @[Top.scala 16:26]
  wire  mmcm_io_CLKOUT1; // @[Top.scala 16:26]
  wire  mmcm_io_CLKIN1_pad_O; // @[Buf.scala 51:34]
  wire  mmcm_io_CLKIN1_pad_I; // @[Buf.scala 51:34]
  wire  mmcm_io_CLKIN1_pad_IB; // @[Buf.scala 51:34]
  wire  hbmDriver_clock; // @[Top.scala 42:71]
  wire  hbmDriver_io_hbm_clk; // @[Top.scala 42:71]
  wire  hbmDriver_io_hbm_rstn; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_aw_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_aw_valid; // @[Top.scala 42:71]
  wire [33:0] hbmDriver_io_axi_hbm_0_aw_bits_addr; // @[Top.scala 42:71]
  wire [3:0] hbmDriver_io_axi_hbm_0_aw_bits_len; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_ar_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_ar_valid; // @[Top.scala 42:71]
  wire [33:0] hbmDriver_io_axi_hbm_0_ar_bits_addr; // @[Top.scala 42:71]
  wire [3:0] hbmDriver_io_axi_hbm_0_ar_bits_len; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_w_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_w_valid; // @[Top.scala 42:71]
  wire [255:0] hbmDriver_io_axi_hbm_0_w_bits_data; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_w_bits_last; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_r_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_0_r_valid; // @[Top.scala 42:71]
  wire [255:0] hbmDriver_io_axi_hbm_0_r_bits_data; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_aw_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_aw_valid; // @[Top.scala 42:71]
  wire [33:0] hbmDriver_io_axi_hbm_1_aw_bits_addr; // @[Top.scala 42:71]
  wire [1:0] hbmDriver_io_axi_hbm_1_aw_bits_burst; // @[Top.scala 42:71]
  wire [3:0] hbmDriver_io_axi_hbm_1_aw_bits_len; // @[Top.scala 42:71]
  wire [2:0] hbmDriver_io_axi_hbm_1_aw_bits_size; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_ar_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_ar_valid; // @[Top.scala 42:71]
  wire [33:0] hbmDriver_io_axi_hbm_1_ar_bits_addr; // @[Top.scala 42:71]
  wire [1:0] hbmDriver_io_axi_hbm_1_ar_bits_burst; // @[Top.scala 42:71]
  wire [3:0] hbmDriver_io_axi_hbm_1_ar_bits_len; // @[Top.scala 42:71]
  wire [2:0] hbmDriver_io_axi_hbm_1_ar_bits_size; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_w_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_w_valid; // @[Top.scala 42:71]
  wire [255:0] hbmDriver_io_axi_hbm_1_w_bits_data; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_w_bits_last; // @[Top.scala 42:71]
  wire [31:0] hbmDriver_io_axi_hbm_1_w_bits_strb; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_r_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_r_valid; // @[Top.scala 42:71]
  wire [255:0] hbmDriver_io_axi_hbm_1_r_bits_data; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_r_bits_last; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_b_ready; // @[Top.scala 42:71]
  wire  hbmDriver_io_axi_hbm_1_b_valid; // @[Top.scala 42:71]
  wire [15:0] qdma_io_pin_tx_p; // @[Top.scala 54:26]
  wire [15:0] qdma_io_pin_tx_n; // @[Top.scala 54:26]
  wire [15:0] qdma_io_pin_rx_p; // @[Top.scala 54:26]
  wire [15:0] qdma_io_pin_rx_n; // @[Top.scala 54:26]
  wire  qdma_io_pin_sys_clk_p; // @[Top.scala 54:26]
  wire  qdma_io_pin_sys_clk_n; // @[Top.scala 54:26]
  wire  qdma_io_pin_sys_rst_n; // @[Top.scala 54:26]
  wire  qdma_io_pcie_clk; // @[Top.scala 54:26]
  wire  qdma_io_pcie_arstn; // @[Top.scala 54:26]
  wire  qdma_io_user_clk; // @[Top.scala 54:26]
  wire  qdma_io_user_arstn; // @[Top.scala 54:26]
  wire  qdma_io_h2c_cmd_ready; // @[Top.scala 54:26]
  wire  qdma_io_h2c_cmd_valid; // @[Top.scala 54:26]
  wire [63:0] qdma_io_h2c_cmd_bits_addr; // @[Top.scala 54:26]
  wire [31:0] qdma_io_h2c_cmd_bits_len; // @[Top.scala 54:26]
  wire  qdma_io_h2c_data_ready; // @[Top.scala 54:26]
  wire  qdma_io_h2c_data_valid; // @[Top.scala 54:26]
  wire [511:0] qdma_io_h2c_data_bits_data; // @[Top.scala 54:26]
  wire  qdma_io_c2h_cmd_ready; // @[Top.scala 54:26]
  wire  qdma_io_c2h_cmd_valid; // @[Top.scala 54:26]
  wire [63:0] qdma_io_c2h_cmd_bits_addr; // @[Top.scala 54:26]
  wire [6:0] qdma_io_c2h_cmd_bits_pfch_tag; // @[Top.scala 54:26]
  wire [31:0] qdma_io_c2h_cmd_bits_len; // @[Top.scala 54:26]
  wire  qdma_io_c2h_data_ready; // @[Top.scala 54:26]
  wire  qdma_io_c2h_data_valid; // @[Top.scala 54:26]
  wire [511:0] qdma_io_c2h_data_bits_data; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_8; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_9; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_10; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_11; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_12; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_13; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_20; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_50; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_51; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_52; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_53; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_54; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_55; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_56; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_57; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_58; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_59; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_70; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_71; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_72; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_73; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_74; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_75; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_76; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_77; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_78; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_79; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_80; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_91; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_92; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_93; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_control_94; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_40; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_51; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_52; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_61; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_71; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_72; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_75; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_76; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_77; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_78; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_79; // @[Top.scala 54:26]
  wire [31:0] qdma_io_reg_status_81; // @[Top.scala 54:26]
  wire  qdma_io_axib_aw_ready; // @[Top.scala 54:26]
  wire  qdma_io_axib_aw_valid; // @[Top.scala 54:26]
  wire [63:0] qdma_io_axib_aw_bits_addr; // @[Top.scala 54:26]
  wire [1:0] qdma_io_axib_aw_bits_burst; // @[Top.scala 54:26]
  wire [7:0] qdma_io_axib_aw_bits_len; // @[Top.scala 54:26]
  wire [2:0] qdma_io_axib_aw_bits_size; // @[Top.scala 54:26]
  wire  qdma_io_axib_ar_ready; // @[Top.scala 54:26]
  wire  qdma_io_axib_ar_valid; // @[Top.scala 54:26]
  wire [63:0] qdma_io_axib_ar_bits_addr; // @[Top.scala 54:26]
  wire [1:0] qdma_io_axib_ar_bits_burst; // @[Top.scala 54:26]
  wire [7:0] qdma_io_axib_ar_bits_len; // @[Top.scala 54:26]
  wire [2:0] qdma_io_axib_ar_bits_size; // @[Top.scala 54:26]
  wire  qdma_io_axib_w_ready; // @[Top.scala 54:26]
  wire  qdma_io_axib_w_valid; // @[Top.scala 54:26]
  wire [511:0] qdma_io_axib_w_bits_data; // @[Top.scala 54:26]
  wire  qdma_io_axib_w_bits_last; // @[Top.scala 54:26]
  wire [63:0] qdma_io_axib_w_bits_strb; // @[Top.scala 54:26]
  wire  qdma_io_axib_r_ready; // @[Top.scala 54:26]
  wire  qdma_io_axib_r_valid; // @[Top.scala 54:26]
  wire [511:0] qdma_io_axib_r_bits_data; // @[Top.scala 54:26]
  wire  qdma_io_axib_r_bits_last; // @[Top.scala 54:26]
  wire  qdma_io_axib_b_valid; // @[Top.scala 54:26]
  wire  qdma_io_c2h_status_last; // @[Top.scala 54:26]
  wire  qdma_io_c2h_status_cmp; // @[Top.scala 54:26]
  wire  qdma_io_c2h_status_valid; // @[Top.scala 54:26]
  wire  qdma_io_c2h_status_error; // @[Top.scala 54:26]
  wire  qdma_io_c2h_status_drop; // @[Top.scala 54:26]
  wire [31:0] qdma_io_tlb_miss_count; // @[Top.scala 54:26]
  wire  h2d_cmd_queue_clock; // @[Top.scala 86:128]
  wire  h2d_cmd_queue_reset; // @[Top.scala 86:128]
  wire  h2d_cmd_queue_io_cmd_in_valid; // @[Top.scala 86:128]
  wire [63:0] h2d_cmd_queue_io_cmd_in_bits_h2c_start_addr; // @[Top.scala 86:128]
  wire [33:0] h2d_cmd_queue_io_cmd_in_bits_h2m_start_addr; // @[Top.scala 86:128]
  wire [31:0] h2d_cmd_queue_io_cmd_in_bits_h2m_length; // @[Top.scala 86:128]
  wire [31:0] h2d_cmd_queue_io_cmd_in_bits_pkt_size; // @[Top.scala 86:128]
  wire [63:0] h2d_cmd_queue_io_cmd_in_bits_h2c_cpt_addr; // @[Top.scala 86:128]
  wire [31:0] h2d_cmd_queue_io_qin; // @[Top.scala 86:128]
  wire  h2d_cmd_queue_io_cmd_out_ready; // @[Top.scala 86:128]
  wire  h2d_cmd_queue_io_cmd_out_valid; // @[Top.scala 86:128]
  wire [63:0] h2d_cmd_queue_io_cmd_out_bits_h2c_start_addr; // @[Top.scala 86:128]
  wire [33:0] h2d_cmd_queue_io_cmd_out_bits_h2m_start_addr; // @[Top.scala 86:128]
  wire [31:0] h2d_cmd_queue_io_cmd_out_bits_h2m_length; // @[Top.scala 86:128]
  wire [63:0] h2d_cmd_queue_io_cmd_out_bits_h2c_cpt_addr; // @[Top.scala 86:128]
  wire [31:0] h2d_cmd_queue_io_h2c_length; // @[Top.scala 86:128]
  wire  h2d_cmd_queue_io_h2m_complete; // @[Top.scala 86:128]
  wire  h2d_cmd_queue_io_h2m_cpt_complete; // @[Top.scala 86:128]
  wire  h2d_cmd_queue_io_last; // @[Top.scala 86:128]
  wire  h2d_cmd_queue_io_h2m_last; // @[Top.scala 86:128]
  wire [31:0] h2d_cmd_queue_io_counter; // @[Top.scala 86:128]
  wire  h2c_clock; // @[Top.scala 98:65]
  wire  h2c_reset; // @[Top.scala 98:65]
  wire [63:0] h2c_io_start_addr; // @[Top.scala 98:65]
  wire [31:0] h2c_io_length; // @[Top.scala 98:65]
  wire  h2c_io_start; // @[Top.scala 98:65]
  wire  h2c_io_h2c_cmd_ready; // @[Top.scala 98:65]
  wire  h2c_io_h2c_cmd_valid; // @[Top.scala 98:65]
  wire [63:0] h2c_io_h2c_cmd_bits_addr; // @[Top.scala 98:65]
  wire [31:0] h2c_io_h2c_cmd_bits_len; // @[Top.scala 98:65]
  wire  h2c_io_complete; // @[Top.scala 98:65]
  wire [31:0] h2c_io_count_time; // @[Top.scala 98:65]
  wire [31:0] h2c_io_send_cmd_count; // @[Top.scala 98:65]
  wire  d2h_cmd_queue_clock; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_reset; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_cmd_in_valid; // @[Top.scala 111:128]
  wire [63:0] d2h_cmd_queue_io_cmd_in_bits_c2h_start_addr; // @[Top.scala 111:128]
  wire [33:0] d2h_cmd_queue_io_cmd_in_bits_m2h_start_addr; // @[Top.scala 111:128]
  wire [31:0] d2h_cmd_queue_io_cmd_in_bits_m2h_length; // @[Top.scala 111:128]
  wire [63:0] d2h_cmd_queue_io_cmd_in_bits_c2h_cpt_addr; // @[Top.scala 111:128]
  wire [31:0] d2h_cmd_queue_io_cmd_in_bits_pkt_size; // @[Top.scala 111:128]
  wire [31:0] d2h_cmd_queue_io_qin; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_cmd_out_ready; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_cmd_out_valid; // @[Top.scala 111:128]
  wire [63:0] d2h_cmd_queue_io_cmd_out_bits_c2h_start_addr; // @[Top.scala 111:128]
  wire [33:0] d2h_cmd_queue_io_cmd_out_bits_m2h_start_addr; // @[Top.scala 111:128]
  wire [31:0] d2h_cmd_queue_io_cmd_out_bits_m2h_length; // @[Top.scala 111:128]
  wire [63:0] d2h_cmd_queue_io_cmd_out_bits_c2h_cpt_addr; // @[Top.scala 111:128]
  wire [31:0] d2h_cmd_queue_io_c2h_length; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_m2h_complete; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_c2h_finish; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_m2h_finish; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_m2h_cpt_complete; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_read_count_equal; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_empty; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_h2m_complete_start; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_h2m_complete; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_h2m_cpt_complete; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_m2h_valid_tmpreg; // @[Top.scala 111:128]
  wire  d2h_cmd_queue_io_last; // @[Top.scala 111:128]
  wire [31:0] d2h_cmd_queue_io_counter; // @[Top.scala 111:128]
  wire  c2h_clock; // @[Top.scala 123:64]
  wire  c2h_reset; // @[Top.scala 123:64]
  wire [63:0] c2h_io_start_addr; // @[Top.scala 123:64]
  wire [31:0] c2h_io_length; // @[Top.scala 123:64]
  wire  c2h_io_start; // @[Top.scala 123:64]
  wire  c2h_io_c2h_cmd_ready; // @[Top.scala 123:64]
  wire  c2h_io_c2h_cmd_valid; // @[Top.scala 123:64]
  wire [63:0] c2h_io_c2h_cmd_bits_addr; // @[Top.scala 123:64]
  wire [6:0] c2h_io_c2h_cmd_bits_pfch_tag; // @[Top.scala 123:64]
  wire [31:0] c2h_io_c2h_cmd_bits_len; // @[Top.scala 123:64]
  wire [31:0] c2h_io_pfch_tag; // @[Top.scala 123:64]
  wire  c2h_io_complete; // @[Top.scala 123:64]
  wire [31:0] c2h_io_count_time; // @[Top.scala 123:64]
  wire [31:0] c2h_io_send_cmd_count; // @[Top.scala 123:64]
  wire  c2h_cpt_clock; // @[Top.scala 137:68]
  wire  c2h_cpt_reset; // @[Top.scala 137:68]
  wire [63:0] c2h_cpt_io_h2c_cpt_addr; // @[Top.scala 137:68]
  wire [63:0] c2h_cpt_io_c2h_cpt_addr; // @[Top.scala 137:68]
  wire [63:0] c2h_cpt_io_p2p_cpt_addr; // @[Top.scala 137:68]
  wire  c2h_cpt_io_h2c_complete; // @[Top.scala 137:68]
  wire  c2h_cpt_io_c2h_complete; // @[Top.scala 137:68]
  wire  c2h_cpt_io_p2p_complete; // @[Top.scala 137:68]
  wire [31:0] c2h_cpt_io_pfch_tag; // @[Top.scala 137:68]
  wire  c2h_cpt_io_h2c_start; // @[Top.scala 137:68]
  wire  c2h_cpt_io_c2h_start; // @[Top.scala 137:68]
  wire  c2h_cpt_io_h2c_cpt_complete; // @[Top.scala 137:68]
  wire  c2h_cpt_io_c2h_cpt_complete; // @[Top.scala 137:68]
  wire  c2h_cpt_io_p2p_cpt_complete; // @[Top.scala 137:68]
  wire [31:0] c2h_cpt_io_polling; // @[Top.scala 137:68]
  wire  c2h_cpt_io_c2h_cmd_ready; // @[Top.scala 137:68]
  wire  c2h_cpt_io_c2h_cmd_valid; // @[Top.scala 137:68]
  wire [63:0] c2h_cpt_io_c2h_cmd_bits_addr; // @[Top.scala 137:68]
  wire [6:0] c2h_cpt_io_c2h_cmd_bits_pfch_tag; // @[Top.scala 137:68]
  wire  c2h_cpt_io_c2h_data_ready; // @[Top.scala 137:68]
  wire  c2h_cpt_io_c2h_data_valid; // @[Top.scala 137:68]
  wire  h2m_clock; // @[Top.scala 165:62]
  wire  h2m_reset; // @[Top.scala 165:62]
  wire [33:0] h2m_io_start_addr; // @[Top.scala 165:62]
  wire [31:0] h2m_io_length; // @[Top.scala 165:62]
  wire  h2m_io_start; // @[Top.scala 165:62]
  wire  h2m_io_complete; // @[Top.scala 165:62]
  wire [33:0] h2m_io_awaddr; // @[Top.scala 165:62]
  wire  h2m_io_awvalid; // @[Top.scala 165:62]
  wire  h2m_io_awready; // @[Top.scala 165:62]
  wire [7:0] h2m_io_awlen; // @[Top.scala 165:62]
  wire  h2m_io_wfire; // @[Top.scala 165:62]
  wire  h2m_io_fifo_rden; // @[Top.scala 165:62]
  wire  h2m_io_wlast; // @[Top.scala 165:62]
  wire  h2m_io_last; // @[Top.scala 165:62]
  wire  h2m_io_clear; // @[Top.scala 165:62]
  wire  m2h_clock; // @[Top.scala 167:62]
  wire  m2h_reset; // @[Top.scala 167:62]
  wire [33:0] m2h_io_start_addr; // @[Top.scala 167:62]
  wire [31:0] m2h_io_length; // @[Top.scala 167:62]
  wire  m2h_io_start; // @[Top.scala 167:62]
  wire  m2h_io_complete; // @[Top.scala 167:62]
  wire [33:0] m2h_io_araddr; // @[Top.scala 167:62]
  wire  m2h_io_arvalid; // @[Top.scala 167:62]
  wire  m2h_io_arready; // @[Top.scala 167:62]
  wire [7:0] m2h_io_arlen; // @[Top.scala 167:62]
  wire  m2h_io_rfire; // @[Top.scala 167:62]
  wire  m2h_io_last; // @[Top.scala 167:62]
  wire  m2h_io_m2h_queue_empty; // @[Top.scala 167:62]
  wire  m2h_io_m2h_valid_tmpreg; // @[Top.scala 167:62]
  wire  m2h_io_read_count_equal; // @[Top.scala 167:62]
  wire [33:0] h2m_start_addr_dest_out; // @[CDC.scala 10:25]
  wire  h2m_start_addr_dest_clk; // @[CDC.scala 10:25]
  wire  h2m_start_addr_src_clk; // @[CDC.scala 10:25]
  wire [33:0] h2m_start_addr_src_in; // @[CDC.scala 10:25]
  wire [31:0] h2m_length_dest_out; // @[CDC.scala 10:25]
  wire  h2m_length_dest_clk; // @[CDC.scala 10:25]
  wire  h2m_length_src_clk; // @[CDC.scala 10:25]
  wire [31:0] h2m_length_src_in; // @[CDC.scala 10:25]
  wire  h2m_last_dest_out; // @[CDC.scala 10:25]
  wire  h2m_last_dest_clk; // @[CDC.scala 10:25]
  wire  h2m_last_src_clk; // @[CDC.scala 10:25]
  wire  h2m_last_src_in; // @[CDC.scala 10:25]
  wire  h2m_start_pulse_dest_pulse; // @[CDC.scala 39:25]
  wire  h2m_start_pulse_dest_clk; // @[CDC.scala 39:25]
  wire  h2m_start_pulse_src_clk; // @[CDC.scala 39:25]
  wire  h2m_start_pulse_src_pulse; // @[CDC.scala 39:25]
  wire  h2m_complete_dest_out; // @[CDC.scala 10:25]
  wire  h2m_complete_dest_clk; // @[CDC.scala 10:25]
  wire  h2m_complete_src_clk; // @[CDC.scala 10:25]
  wire  h2m_complete_src_in; // @[CDC.scala 10:25]
  wire  h2m_clear_dest_out; // @[CDC.scala 10:25]
  wire  h2m_clear_dest_clk; // @[CDC.scala 10:25]
  wire  h2m_clear_src_clk; // @[CDC.scala 10:25]
  wire  h2m_clear_src_in; // @[CDC.scala 10:25]
  wire  h2m_cmd_buffer_clock; // @[XQueue.scala 35:23]
  wire  h2m_cmd_buffer_reset; // @[XQueue.scala 35:23]
  wire  h2m_cmd_buffer_io_in_ready; // @[XQueue.scala 35:23]
  wire  h2m_cmd_buffer_io_in_valid; // @[XQueue.scala 35:23]
  wire [66:0] h2m_cmd_buffer_io_in_bits; // @[XQueue.scala 35:23]
  wire  h2m_cmd_buffer_io_out_ready; // @[XQueue.scala 35:23]
  wire  h2m_cmd_buffer_io_out_valid; // @[XQueue.scala 35:23]
  wire [66:0] h2m_cmd_buffer_io_out_bits; // @[XQueue.scala 35:23]
  wire  h2m_cmd_buffer_ready_clock; // @[Top.scala 184:120]
  wire  h2m_cmd_buffer_ready_reset; // @[Top.scala 184:120]
  wire  h2m_cmd_buffer_ready_io_ready; // @[Top.scala 184:120]
  wire  h2m_cmd_buffer_ready_io_valid; // @[Top.scala 184:120]
  wire  h2m_cmd_buffer_ready_io_complete; // @[Top.scala 184:120]
  wire [63:0] m2h_start_addr_dest_out; // @[CDC.scala 10:25]
  wire  m2h_start_addr_dest_clk; // @[CDC.scala 10:25]
  wire  m2h_start_addr_src_clk; // @[CDC.scala 10:25]
  wire [63:0] m2h_start_addr_src_in; // @[CDC.scala 10:25]
  wire [31:0] m2h_length_dest_out; // @[CDC.scala 10:25]
  wire  m2h_length_dest_clk; // @[CDC.scala 10:25]
  wire  m2h_length_src_clk; // @[CDC.scala 10:25]
  wire [31:0] m2h_length_src_in; // @[CDC.scala 10:25]
  wire  m2h_start_pulse_dest_pulse; // @[CDC.scala 39:25]
  wire  m2h_start_pulse_dest_clk; // @[CDC.scala 39:25]
  wire  m2h_start_pulse_src_clk; // @[CDC.scala 39:25]
  wire  m2h_start_pulse_src_pulse; // @[CDC.scala 39:25]
  wire  m2h_complete_dest_out; // @[CDC.scala 10:25]
  wire  m2h_complete_dest_clk; // @[CDC.scala 10:25]
  wire  m2h_complete_src_clk; // @[CDC.scala 10:25]
  wire  m2h_complete_src_in; // @[CDC.scala 10:25]
  wire  m2h_last_dest_out; // @[CDC.scala 10:25]
  wire  m2h_last_dest_clk; // @[CDC.scala 10:25]
  wire  m2h_last_src_clk; // @[CDC.scala 10:25]
  wire  m2h_last_src_in; // @[CDC.scala 10:25]
  wire  m2h_read_count_equal_dest_out; // @[CDC.scala 10:25]
  wire  m2h_read_count_equal_dest_clk; // @[CDC.scala 10:25]
  wire  m2h_read_count_equal_src_clk; // @[CDC.scala 10:25]
  wire  m2h_read_count_equal_src_in; // @[CDC.scala 10:25]
  wire  c2h_status_clock; // @[Top.scala 244:129]
  wire  c2h_status_reset; // @[Top.scala 244:129]
  wire  c2h_status_io_c2h_start; // @[Top.scala 244:129]
  wire  c2h_status_io_c2h_status_last; // @[Top.scala 244:129]
  wire  c2h_status_io_c2h_status_cmp; // @[Top.scala 244:129]
  wire  c2h_status_io_c2h_status_valid; // @[Top.scala 244:129]
  wire  c2h_status_io_c2h_status_error; // @[Top.scala 244:129]
  wire  c2h_status_io_c2h_status_drop; // @[Top.scala 244:129]
  wire [31:0] c2h_status_io_c2h_status_last_count; // @[Top.scala 244:129]
  wire [31:0] c2h_status_io_c2h_status_cmp_count; // @[Top.scala 244:129]
  wire [31:0] c2h_status_io_c2h_status_valid_count; // @[Top.scala 244:129]
  wire [31:0] c2h_status_io_c2h_status_error_count; // @[Top.scala 244:129]
  wire [31:0] c2h_status_io_c2h_status_drop_count; // @[Top.scala 244:129]
  wire  c2h_status_start_dest_out; // @[CDC.scala 10:25]
  wire  c2h_status_start_dest_clk; // @[CDC.scala 10:25]
  wire  c2h_status_start_src_clk; // @[CDC.scala 10:25]
  wire  c2h_status_start_src_in; // @[CDC.scala 10:25]
  wire [31:0] last_count_dest_out; // @[CDC.scala 10:25]
  wire  last_count_dest_clk; // @[CDC.scala 10:25]
  wire  last_count_src_clk; // @[CDC.scala 10:25]
  wire [31:0] last_count_src_in; // @[CDC.scala 10:25]
  wire [31:0] cmp_count_dest_out; // @[CDC.scala 10:25]
  wire  cmp_count_dest_clk; // @[CDC.scala 10:25]
  wire  cmp_count_src_clk; // @[CDC.scala 10:25]
  wire [31:0] cmp_count_src_in; // @[CDC.scala 10:25]
  wire [31:0] valid_count_dest_out; // @[CDC.scala 10:25]
  wire  valid_count_dest_clk; // @[CDC.scala 10:25]
  wire  valid_count_src_clk; // @[CDC.scala 10:25]
  wire [31:0] valid_count_src_in; // @[CDC.scala 10:25]
  wire [31:0] error_count_dest_out; // @[CDC.scala 10:25]
  wire  error_count_dest_clk; // @[CDC.scala 10:25]
  wire  error_count_src_clk; // @[CDC.scala 10:25]
  wire [31:0] error_count_src_in; // @[CDC.scala 10:25]
  wire [31:0] drop_count_dest_out; // @[CDC.scala 10:25]
  wire  drop_count_dest_clk; // @[CDC.scala 10:25]
  wire  drop_count_src_clk; // @[CDC.scala 10:25]
  wire [31:0] drop_count_src_in; // @[CDC.scala 10:25]
  wire  h2m_queue_almost_empty; // @[Top.scala 275:31]
  wire  h2m_queue_almost_full; // @[Top.scala 275:31]
  wire  h2m_queue_data_valid; // @[Top.scala 275:31]
  wire  h2m_queue_dbiterr; // @[Top.scala 275:31]
  wire [255:0] h2m_queue_dout; // @[Top.scala 275:31]
  wire  h2m_queue_empty; // @[Top.scala 275:31]
  wire  h2m_queue_full; // @[Top.scala 275:31]
  wire  h2m_queue_overflow; // @[Top.scala 275:31]
  wire  h2m_queue_prog_empty; // @[Top.scala 275:31]
  wire  h2m_queue_prog_full; // @[Top.scala 275:31]
  wire  h2m_queue_rd_data_count; // @[Top.scala 275:31]
  wire  h2m_queue_rd_rst_busy; // @[Top.scala 275:31]
  wire  h2m_queue_sbiterr; // @[Top.scala 275:31]
  wire  h2m_queue_underflow; // @[Top.scala 275:31]
  wire  h2m_queue_wr_ack; // @[Top.scala 275:31]
  wire  h2m_queue_wr_data_count; // @[Top.scala 275:31]
  wire  h2m_queue_wr_rst_busy; // @[Top.scala 275:31]
  wire [511:0] h2m_queue_din; // @[Top.scala 275:31]
  wire  h2m_queue_injectdbiterr; // @[Top.scala 275:31]
  wire  h2m_queue_injectsbiterr; // @[Top.scala 275:31]
  wire  h2m_queue_rd_clk; // @[Top.scala 275:31]
  wire  h2m_queue_rd_en; // @[Top.scala 275:31]
  wire  h2m_queue_rst; // @[Top.scala 275:31]
  wire  h2m_queue_sleep; // @[Top.scala 275:31]
  wire  h2m_queue_wr_clk; // @[Top.scala 275:31]
  wire  h2m_queue_wr_en; // @[Top.scala 275:31]
  wire  m2h_queue__almost_empty; // @[Top.scala 276:31]
  wire  m2h_queue__almost_full; // @[Top.scala 276:31]
  wire  m2h_queue__data_valid; // @[Top.scala 276:31]
  wire  m2h_queue__dbiterr; // @[Top.scala 276:31]
  wire [511:0] m2h_queue__dout; // @[Top.scala 276:31]
  wire  m2h_queue__empty; // @[Top.scala 276:31]
  wire  m2h_queue__full; // @[Top.scala 276:31]
  wire  m2h_queue__overflow; // @[Top.scala 276:31]
  wire  m2h_queue__prog_empty; // @[Top.scala 276:31]
  wire  m2h_queue__prog_full; // @[Top.scala 276:31]
  wire  m2h_queue__rd_data_count; // @[Top.scala 276:31]
  wire  m2h_queue__rd_rst_busy; // @[Top.scala 276:31]
  wire  m2h_queue__sbiterr; // @[Top.scala 276:31]
  wire  m2h_queue__underflow; // @[Top.scala 276:31]
  wire  m2h_queue__wr_ack; // @[Top.scala 276:31]
  wire  m2h_queue__wr_data_count; // @[Top.scala 276:31]
  wire  m2h_queue__wr_rst_busy; // @[Top.scala 276:31]
  wire [255:0] m2h_queue__din; // @[Top.scala 276:31]
  wire  m2h_queue__injectdbiterr; // @[Top.scala 276:31]
  wire  m2h_queue__injectsbiterr; // @[Top.scala 276:31]
  wire  m2h_queue__rd_clk; // @[Top.scala 276:31]
  wire  m2h_queue__rd_en; // @[Top.scala 276:31]
  wire  m2h_queue__rst; // @[Top.scala 276:31]
  wire  m2h_queue__sleep; // @[Top.scala 276:31]
  wire  m2h_queue__wr_clk; // @[Top.scala 276:31]
  wire  m2h_queue__wr_en; // @[Top.scala 276:31]
  wire  h2m_valid_tmpreg_clock; // @[Top.scala 289:118]
  wire  h2m_valid_tmpreg_reset; // @[Top.scala 289:118]
  wire  h2m_valid_tmpreg_io_ready; // @[Top.scala 289:118]
  wire  h2m_valid_tmpreg_io_valid; // @[Top.scala 289:118]
  wire  h2m_valid_tmpreg_io_tmpreg; // @[Top.scala 289:118]
  wire  m2h_valid_tmpreg_clock; // @[Top.scala 305:120]
  wire  m2h_valid_tmpreg_reset; // @[Top.scala 305:120]
  wire  m2h_valid_tmpreg_io_ready; // @[Top.scala 305:120]
  wire  m2h_valid_tmpreg_io_valid; // @[Top.scala 305:120]
  wire  m2h_valid_tmpreg_io_tmpreg; // @[Top.scala 305:120]
  wire  m2h_queue_empty_dest_out; // @[CDC.scala 10:25]
  wire  m2h_queue_empty_dest_clk; // @[CDC.scala 10:25]
  wire  m2h_queue_empty_src_clk; // @[CDC.scala 10:25]
  wire  m2h_queue_empty_src_in; // @[CDC.scala 10:25]
  wire  m2h_valid_tmpreg_tom2h_dest_out; // @[CDC.scala 10:25]
  wire  m2h_valid_tmpreg_tom2h_dest_clk; // @[CDC.scala 10:25]
  wire  m2h_valid_tmpreg_tom2h_src_clk; // @[CDC.scala 10:25]
  wire  m2h_valid_tmpreg_tom2h_src_in; // @[CDC.scala 10:25]
  wire [63:0] axicc_s_axi_awaddr; // @[Top.scala 356:27]
  wire [7:0] axicc_s_axi_awlen; // @[Top.scala 356:27]
  wire [2:0] axicc_s_axi_awsize; // @[Top.scala 356:27]
  wire [1:0] axicc_s_axi_awburst; // @[Top.scala 356:27]
  wire  axicc_s_axi_awlock; // @[Top.scala 356:27]
  wire [3:0] axicc_s_axi_awcache; // @[Top.scala 356:27]
  wire [2:0] axicc_s_axi_awprot; // @[Top.scala 356:27]
  wire [3:0] axicc_s_axi_awregion; // @[Top.scala 356:27]
  wire [3:0] axicc_s_axi_awqos; // @[Top.scala 356:27]
  wire  axicc_s_axi_awvalid; // @[Top.scala 356:27]
  wire  axicc_s_axi_awready; // @[Top.scala 356:27]
  wire [511:0] axicc_s_axi_wdata; // @[Top.scala 356:27]
  wire [63:0] axicc_s_axi_wstrb; // @[Top.scala 356:27]
  wire  axicc_s_axi_wlast; // @[Top.scala 356:27]
  wire  axicc_s_axi_wvalid; // @[Top.scala 356:27]
  wire  axicc_s_axi_wready; // @[Top.scala 356:27]
  wire [1:0] axicc_s_axi_bresp; // @[Top.scala 356:27]
  wire  axicc_s_axi_bvalid; // @[Top.scala 356:27]
  wire  axicc_s_axi_bready; // @[Top.scala 356:27]
  wire [63:0] axicc_s_axi_araddr; // @[Top.scala 356:27]
  wire [7:0] axicc_s_axi_arlen; // @[Top.scala 356:27]
  wire [2:0] axicc_s_axi_arsize; // @[Top.scala 356:27]
  wire [1:0] axicc_s_axi_arburst; // @[Top.scala 356:27]
  wire  axicc_s_axi_arlock; // @[Top.scala 356:27]
  wire [3:0] axicc_s_axi_arcache; // @[Top.scala 356:27]
  wire [2:0] axicc_s_axi_arprot; // @[Top.scala 356:27]
  wire [3:0] axicc_s_axi_arregion; // @[Top.scala 356:27]
  wire [3:0] axicc_s_axi_arqos; // @[Top.scala 356:27]
  wire  axicc_s_axi_arvalid; // @[Top.scala 356:27]
  wire  axicc_s_axi_arready; // @[Top.scala 356:27]
  wire [511:0] axicc_s_axi_rdata; // @[Top.scala 356:27]
  wire [1:0] axicc_s_axi_rresp; // @[Top.scala 356:27]
  wire  axicc_s_axi_rlast; // @[Top.scala 356:27]
  wire  axicc_s_axi_rvalid; // @[Top.scala 356:27]
  wire  axicc_s_axi_rready; // @[Top.scala 356:27]
  wire  axicc_s_axi_aclk; // @[Top.scala 356:27]
  wire  axicc_s_axi_aresetn; // @[Top.scala 356:27]
  wire  axicc_m_axi_aclk; // @[Top.scala 356:27]
  wire  axicc_m_axi_aresetn; // @[Top.scala 356:27]
  wire [63:0] axicc_m_axi_awaddr; // @[Top.scala 356:27]
  wire [7:0] axicc_m_axi_awlen; // @[Top.scala 356:27]
  wire [2:0] axicc_m_axi_awsize; // @[Top.scala 356:27]
  wire [1:0] axicc_m_axi_awburst; // @[Top.scala 356:27]
  wire  axicc_m_axi_awlock; // @[Top.scala 356:27]
  wire [3:0] axicc_m_axi_awcache; // @[Top.scala 356:27]
  wire [2:0] axicc_m_axi_awprot; // @[Top.scala 356:27]
  wire [3:0] axicc_m_axi_awregion; // @[Top.scala 356:27]
  wire [3:0] axicc_m_axi_awqos; // @[Top.scala 356:27]
  wire  axicc_m_axi_awvalid; // @[Top.scala 356:27]
  wire  axicc_m_axi_awready; // @[Top.scala 356:27]
  wire [511:0] axicc_m_axi_wdata; // @[Top.scala 356:27]
  wire [63:0] axicc_m_axi_wstrb; // @[Top.scala 356:27]
  wire  axicc_m_axi_wlast; // @[Top.scala 356:27]
  wire  axicc_m_axi_wvalid; // @[Top.scala 356:27]
  wire  axicc_m_axi_wready; // @[Top.scala 356:27]
  wire [1:0] axicc_m_axi_bresp; // @[Top.scala 356:27]
  wire  axicc_m_axi_bvalid; // @[Top.scala 356:27]
  wire  axicc_m_axi_bready; // @[Top.scala 356:27]
  wire [63:0] axicc_m_axi_araddr; // @[Top.scala 356:27]
  wire [7:0] axicc_m_axi_arlen; // @[Top.scala 356:27]
  wire [2:0] axicc_m_axi_arsize; // @[Top.scala 356:27]
  wire [1:0] axicc_m_axi_arburst; // @[Top.scala 356:27]
  wire  axicc_m_axi_arlock; // @[Top.scala 356:27]
  wire [3:0] axicc_m_axi_arcache; // @[Top.scala 356:27]
  wire [2:0] axicc_m_axi_arprot; // @[Top.scala 356:27]
  wire [3:0] axicc_m_axi_arregion; // @[Top.scala 356:27]
  wire [3:0] axicc_m_axi_arqos; // @[Top.scala 356:27]
  wire  axicc_m_axi_arvalid; // @[Top.scala 356:27]
  wire  axicc_m_axi_arready; // @[Top.scala 356:27]
  wire [511:0] axicc_m_axi_rdata; // @[Top.scala 356:27]
  wire [1:0] axicc_m_axi_rresp; // @[Top.scala 356:27]
  wire  axicc_m_axi_rlast; // @[Top.scala 356:27]
  wire  axicc_m_axi_rvalid; // @[Top.scala 356:27]
  wire  axicc_m_axi_rready; // @[Top.scala 356:27]
  wire [33:0] axidwc_s_axi_awaddr; // @[Top.scala 404:28]
  wire [7:0] axidwc_s_axi_awlen; // @[Top.scala 404:28]
  wire [2:0] axidwc_s_axi_awsize; // @[Top.scala 404:28]
  wire [1:0] axidwc_s_axi_awburst; // @[Top.scala 404:28]
  wire  axidwc_s_axi_awlock; // @[Top.scala 404:28]
  wire [3:0] axidwc_s_axi_awcache; // @[Top.scala 404:28]
  wire [2:0] axidwc_s_axi_awprot; // @[Top.scala 404:28]
  wire [3:0] axidwc_s_axi_awregion; // @[Top.scala 404:28]
  wire [3:0] axidwc_s_axi_awqos; // @[Top.scala 404:28]
  wire  axidwc_s_axi_awvalid; // @[Top.scala 404:28]
  wire  axidwc_s_axi_awready; // @[Top.scala 404:28]
  wire [511:0] axidwc_s_axi_wdata; // @[Top.scala 404:28]
  wire [63:0] axidwc_s_axi_wstrb; // @[Top.scala 404:28]
  wire  axidwc_s_axi_wlast; // @[Top.scala 404:28]
  wire  axidwc_s_axi_wvalid; // @[Top.scala 404:28]
  wire  axidwc_s_axi_wready; // @[Top.scala 404:28]
  wire [1:0] axidwc_s_axi_bresp; // @[Top.scala 404:28]
  wire  axidwc_s_axi_bvalid; // @[Top.scala 404:28]
  wire  axidwc_s_axi_bready; // @[Top.scala 404:28]
  wire [33:0] axidwc_s_axi_araddr; // @[Top.scala 404:28]
  wire [7:0] axidwc_s_axi_arlen; // @[Top.scala 404:28]
  wire [2:0] axidwc_s_axi_arsize; // @[Top.scala 404:28]
  wire [1:0] axidwc_s_axi_arburst; // @[Top.scala 404:28]
  wire  axidwc_s_axi_arlock; // @[Top.scala 404:28]
  wire [3:0] axidwc_s_axi_arcache; // @[Top.scala 404:28]
  wire [2:0] axidwc_s_axi_arprot; // @[Top.scala 404:28]
  wire [3:0] axidwc_s_axi_arregion; // @[Top.scala 404:28]
  wire [3:0] axidwc_s_axi_arqos; // @[Top.scala 404:28]
  wire  axidwc_s_axi_arvalid; // @[Top.scala 404:28]
  wire  axidwc_s_axi_arready; // @[Top.scala 404:28]
  wire [511:0] axidwc_s_axi_rdata; // @[Top.scala 404:28]
  wire [1:0] axidwc_s_axi_rresp; // @[Top.scala 404:28]
  wire  axidwc_s_axi_rlast; // @[Top.scala 404:28]
  wire  axidwc_s_axi_rvalid; // @[Top.scala 404:28]
  wire  axidwc_s_axi_rready; // @[Top.scala 404:28]
  wire  axidwc_s_axi_aclk; // @[Top.scala 404:28]
  wire  axidwc_s_axi_aresetn; // @[Top.scala 404:28]
  wire [33:0] axidwc_m_axi_awaddr; // @[Top.scala 404:28]
  wire [7:0] axidwc_m_axi_awlen; // @[Top.scala 404:28]
  wire [2:0] axidwc_m_axi_awsize; // @[Top.scala 404:28]
  wire [1:0] axidwc_m_axi_awburst; // @[Top.scala 404:28]
  wire  axidwc_m_axi_awlock; // @[Top.scala 404:28]
  wire [3:0] axidwc_m_axi_awcache; // @[Top.scala 404:28]
  wire [2:0] axidwc_m_axi_awprot; // @[Top.scala 404:28]
  wire [3:0] axidwc_m_axi_awregion; // @[Top.scala 404:28]
  wire [3:0] axidwc_m_axi_awqos; // @[Top.scala 404:28]
  wire  axidwc_m_axi_awvalid; // @[Top.scala 404:28]
  wire  axidwc_m_axi_awready; // @[Top.scala 404:28]
  wire [255:0] axidwc_m_axi_wdata; // @[Top.scala 404:28]
  wire [31:0] axidwc_m_axi_wstrb; // @[Top.scala 404:28]
  wire  axidwc_m_axi_wlast; // @[Top.scala 404:28]
  wire  axidwc_m_axi_wvalid; // @[Top.scala 404:28]
  wire  axidwc_m_axi_wready; // @[Top.scala 404:28]
  wire [1:0] axidwc_m_axi_bresp; // @[Top.scala 404:28]
  wire  axidwc_m_axi_bvalid; // @[Top.scala 404:28]
  wire  axidwc_m_axi_bready; // @[Top.scala 404:28]
  wire [33:0] axidwc_m_axi_araddr; // @[Top.scala 404:28]
  wire [7:0] axidwc_m_axi_arlen; // @[Top.scala 404:28]
  wire [2:0] axidwc_m_axi_arsize; // @[Top.scala 404:28]
  wire [1:0] axidwc_m_axi_arburst; // @[Top.scala 404:28]
  wire  axidwc_m_axi_arlock; // @[Top.scala 404:28]
  wire [3:0] axidwc_m_axi_arcache; // @[Top.scala 404:28]
  wire [2:0] axidwc_m_axi_arprot; // @[Top.scala 404:28]
  wire [3:0] axidwc_m_axi_arregion; // @[Top.scala 404:28]
  wire [3:0] axidwc_m_axi_arqos; // @[Top.scala 404:28]
  wire  axidwc_m_axi_arvalid; // @[Top.scala 404:28]
  wire  axidwc_m_axi_arready; // @[Top.scala 404:28]
  wire [255:0] axidwc_m_axi_rdata; // @[Top.scala 404:28]
  wire [1:0] axidwc_m_axi_rresp; // @[Top.scala 404:28]
  wire  axidwc_m_axi_rlast; // @[Top.scala 404:28]
  wire  axidwc_m_axi_rvalid; // @[Top.scala 404:28]
  wire  axidwc_m_axi_rready; // @[Top.scala 404:28]
  wire  p2p_counter_clock; // @[Top.scala 472:102]
  wire  p2p_counter_reset; // @[Top.scala 472:102]
  wire  p2p_counter_io_start; // @[Top.scala 472:102]
  wire [31:0] p2p_counter_io_length; // @[Top.scala 472:102]
  wire  p2p_counter_io_wready; // @[Top.scala 472:102]
  wire  p2p_counter_io_wvalid; // @[Top.scala 472:102]
  wire [31:0] p2p_counter_io_wdatasample; // @[Top.scala 472:102]
  wire  p2p_counter_io_p2p_complete; // @[Top.scala 472:102]
  wire  p2p_counter_io_p2p_cpt_complete; // @[Top.scala 472:102]
  wire [63:0] p2p_cpt_addr_dest_out; // @[CDC.scala 10:25]
  wire  p2p_cpt_addr_dest_clk; // @[CDC.scala 10:25]
  wire  p2p_cpt_addr_src_clk; // @[CDC.scala 10:25]
  wire [63:0] p2p_cpt_addr_src_in; // @[CDC.scala 10:25]
  wire [31:0] p2p_length_dest_out; // @[CDC.scala 10:25]
  wire  p2p_length_dest_clk; // @[CDC.scala 10:25]
  wire  p2p_length_src_clk; // @[CDC.scala 10:25]
  wire [31:0] p2p_length_src_in; // @[CDC.scala 10:25]
  wire  p2p_start_dest_out; // @[CDC.scala 10:25]
  wire  p2p_start_dest_clk; // @[CDC.scala 10:25]
  wire  p2p_start_src_clk; // @[CDC.scala 10:25]
  wire  p2p_start_src_in; // @[CDC.scala 10:25]
  wire  p2p_complete_dest_pulse; // @[CDC.scala 39:25]
  wire  p2p_complete_dest_clk; // @[CDC.scala 39:25]
  wire  p2p_complete_src_clk; // @[CDC.scala 39:25]
  wire  p2p_complete_src_pulse; // @[CDC.scala 39:25]
  wire  p2p_cpt_complete_dest_pulse; // @[CDC.scala 39:25]
  wire  p2p_cpt_complete_dest_clk; // @[CDC.scala 39:25]
  wire  p2p_cpt_complete_src_clk; // @[CDC.scala 39:25]
  wire  p2p_cpt_complete_src_pulse; // @[CDC.scala 39:25]
  reg  hbm_rstn; // @[Top.scala 45:70]
  wire  _T = ~mmcm_io_LOCKED; // @[Top.scala 86:110]
  reg  h2d_cmd_queue_io_cmd_in_valid_REG; // @[Top.scala 95:141]
  reg  h2d_cmd_queue_io_cmd_in_valid_REG_1; // @[Top.scala 95:133]
  reg  h2d_cmd_queue_io_cmd_in_valid_REG_2; // @[Top.scala 95:125]
  reg  h2d_cmd_queue_io_cmd_in_valid_REG_3; // @[Top.scala 37:48]
  reg  d2h_cmd_queue_io_cmd_in_valid_REG; // @[Top.scala 120:141]
  reg  d2h_cmd_queue_io_cmd_in_valid_REG_1; // @[Top.scala 120:133]
  reg  d2h_cmd_queue_io_cmd_in_valid_REG_2; // @[Top.scala 120:125]
  reg  d2h_cmd_queue_io_cmd_in_valid_REG_3; // @[Top.scala 37:48]
  reg  c2h_cpt_io_h2c_start_REG; // @[Top.scala 37:48]
  reg  c2h_cpt_io_c2h_start_REG; // @[Top.scala 37:48]
  reg  d2h_cmd_queue_io_h2m_complete_start_REG; // @[Top.scala 37:48]
  wire  _c2h_io_c2h_cmd_ready_T = ~c2h_cpt_io_c2h_cmd_valid; // @[Top.scala 157:100]
  wire [34:0] h2m_cmd_buffer_io_in_bits_hi = {h2d_cmd_queue_io_h2m_last,h2d_cmd_queue_io_cmd_out_bits_h2m_start_addr}; // @[Cat.scala 30:58]
  reg [33:0] h2m_start_addr_reg; // @[Top.scala 189:121]
  reg [33:0] h2m_length_reg; // @[Top.scala 190:129]
  reg  h2m_last_reg; // @[Top.scala 191:129]
  wire  _T_9 = h2m_cmd_buffer_io_out_ready & h2m_cmd_buffer_io_out_valid; // @[Decoupled.scala 40:37]
  reg  h2m_io_start_REG; // @[Top.scala 206:128]
  reg  m2h_io_start_REG; // @[Top.scala 224:128]
  wire  pcie_rstn = qdma_io_pcie_arstn; // @[Top.scala 64:39 Top.scala 66:41]
  reg  p2p_start_io_src_in_REG; // @[Top.scala 484:115]
  reg  p2p_start_io_src_in_REG_1; // @[Top.scala 484:107]
  reg  p2p_start_io_src_in_REG_2; // @[Top.scala 484:99]
  reg  p2p_counter_io_start_REG; // @[Top.scala 485:96]
  MMCME4_ADV_Wrapper mmcm ( // @[Top.scala 16:26]
    .io_CLKIN1(mmcm_io_CLKIN1),
    .io_LOCKED(mmcm_io_LOCKED),
    .io_CLKOUT0(mmcm_io_CLKOUT0),
    .io_CLKOUT1(mmcm_io_CLKOUT1)
  );
  IBUFDS mmcm_io_CLKIN1_pad ( // @[Buf.scala 51:34]
    .O(mmcm_io_CLKIN1_pad_O),
    .I(mmcm_io_CLKIN1_pad_I),
    .IB(mmcm_io_CLKIN1_pad_IB)
  );
  HBM_DRIVER hbmDriver ( // @[Top.scala 42:71]
    .clock(hbmDriver_clock),
    .io_hbm_clk(hbmDriver_io_hbm_clk),
    .io_hbm_rstn(hbmDriver_io_hbm_rstn),
    .io_axi_hbm_0_aw_ready(hbmDriver_io_axi_hbm_0_aw_ready),
    .io_axi_hbm_0_aw_valid(hbmDriver_io_axi_hbm_0_aw_valid),
    .io_axi_hbm_0_aw_bits_addr(hbmDriver_io_axi_hbm_0_aw_bits_addr),
    .io_axi_hbm_0_aw_bits_len(hbmDriver_io_axi_hbm_0_aw_bits_len),
    .io_axi_hbm_0_ar_ready(hbmDriver_io_axi_hbm_0_ar_ready),
    .io_axi_hbm_0_ar_valid(hbmDriver_io_axi_hbm_0_ar_valid),
    .io_axi_hbm_0_ar_bits_addr(hbmDriver_io_axi_hbm_0_ar_bits_addr),
    .io_axi_hbm_0_ar_bits_len(hbmDriver_io_axi_hbm_0_ar_bits_len),
    .io_axi_hbm_0_w_ready(hbmDriver_io_axi_hbm_0_w_ready),
    .io_axi_hbm_0_w_valid(hbmDriver_io_axi_hbm_0_w_valid),
    .io_axi_hbm_0_w_bits_data(hbmDriver_io_axi_hbm_0_w_bits_data),
    .io_axi_hbm_0_w_bits_last(hbmDriver_io_axi_hbm_0_w_bits_last),
    .io_axi_hbm_0_r_ready(hbmDriver_io_axi_hbm_0_r_ready),
    .io_axi_hbm_0_r_valid(hbmDriver_io_axi_hbm_0_r_valid),
    .io_axi_hbm_0_r_bits_data(hbmDriver_io_axi_hbm_0_r_bits_data),
    .io_axi_hbm_1_aw_ready(hbmDriver_io_axi_hbm_1_aw_ready),
    .io_axi_hbm_1_aw_valid(hbmDriver_io_axi_hbm_1_aw_valid),
    .io_axi_hbm_1_aw_bits_addr(hbmDriver_io_axi_hbm_1_aw_bits_addr),
    .io_axi_hbm_1_aw_bits_burst(hbmDriver_io_axi_hbm_1_aw_bits_burst),
    .io_axi_hbm_1_aw_bits_len(hbmDriver_io_axi_hbm_1_aw_bits_len),
    .io_axi_hbm_1_aw_bits_size(hbmDriver_io_axi_hbm_1_aw_bits_size),
    .io_axi_hbm_1_ar_ready(hbmDriver_io_axi_hbm_1_ar_ready),
    .io_axi_hbm_1_ar_valid(hbmDriver_io_axi_hbm_1_ar_valid),
    .io_axi_hbm_1_ar_bits_addr(hbmDriver_io_axi_hbm_1_ar_bits_addr),
    .io_axi_hbm_1_ar_bits_burst(hbmDriver_io_axi_hbm_1_ar_bits_burst),
    .io_axi_hbm_1_ar_bits_len(hbmDriver_io_axi_hbm_1_ar_bits_len),
    .io_axi_hbm_1_ar_bits_size(hbmDriver_io_axi_hbm_1_ar_bits_size),
    .io_axi_hbm_1_w_ready(hbmDriver_io_axi_hbm_1_w_ready),
    .io_axi_hbm_1_w_valid(hbmDriver_io_axi_hbm_1_w_valid),
    .io_axi_hbm_1_w_bits_data(hbmDriver_io_axi_hbm_1_w_bits_data),
    .io_axi_hbm_1_w_bits_last(hbmDriver_io_axi_hbm_1_w_bits_last),
    .io_axi_hbm_1_w_bits_strb(hbmDriver_io_axi_hbm_1_w_bits_strb),
    .io_axi_hbm_1_r_ready(hbmDriver_io_axi_hbm_1_r_ready),
    .io_axi_hbm_1_r_valid(hbmDriver_io_axi_hbm_1_r_valid),
    .io_axi_hbm_1_r_bits_data(hbmDriver_io_axi_hbm_1_r_bits_data),
    .io_axi_hbm_1_r_bits_last(hbmDriver_io_axi_hbm_1_r_bits_last),
    .io_axi_hbm_1_b_ready(hbmDriver_io_axi_hbm_1_b_ready),
    .io_axi_hbm_1_b_valid(hbmDriver_io_axi_hbm_1_b_valid)
  );
  QDMA qdma ( // @[Top.scala 54:26]
    .io_pin_tx_p(qdma_io_pin_tx_p),
    .io_pin_tx_n(qdma_io_pin_tx_n),
    .io_pin_rx_p(qdma_io_pin_rx_p),
    .io_pin_rx_n(qdma_io_pin_rx_n),
    .io_pin_sys_clk_p(qdma_io_pin_sys_clk_p),
    .io_pin_sys_clk_n(qdma_io_pin_sys_clk_n),
    .io_pin_sys_rst_n(qdma_io_pin_sys_rst_n),
    .io_pcie_clk(qdma_io_pcie_clk),
    .io_pcie_arstn(qdma_io_pcie_arstn),
    .io_user_clk(qdma_io_user_clk),
    .io_user_arstn(qdma_io_user_arstn),
    .io_h2c_cmd_ready(qdma_io_h2c_cmd_ready),
    .io_h2c_cmd_valid(qdma_io_h2c_cmd_valid),
    .io_h2c_cmd_bits_addr(qdma_io_h2c_cmd_bits_addr),
    .io_h2c_cmd_bits_len(qdma_io_h2c_cmd_bits_len),
    .io_h2c_data_ready(qdma_io_h2c_data_ready),
    .io_h2c_data_valid(qdma_io_h2c_data_valid),
    .io_h2c_data_bits_data(qdma_io_h2c_data_bits_data),
    .io_c2h_cmd_ready(qdma_io_c2h_cmd_ready),
    .io_c2h_cmd_valid(qdma_io_c2h_cmd_valid),
    .io_c2h_cmd_bits_addr(qdma_io_c2h_cmd_bits_addr),
    .io_c2h_cmd_bits_pfch_tag(qdma_io_c2h_cmd_bits_pfch_tag),
    .io_c2h_cmd_bits_len(qdma_io_c2h_cmd_bits_len),
    .io_c2h_data_ready(qdma_io_c2h_data_ready),
    .io_c2h_data_valid(qdma_io_c2h_data_valid),
    .io_c2h_data_bits_data(qdma_io_c2h_data_bits_data),
    .io_reg_control_8(qdma_io_reg_control_8),
    .io_reg_control_9(qdma_io_reg_control_9),
    .io_reg_control_10(qdma_io_reg_control_10),
    .io_reg_control_11(qdma_io_reg_control_11),
    .io_reg_control_12(qdma_io_reg_control_12),
    .io_reg_control_13(qdma_io_reg_control_13),
    .io_reg_control_20(qdma_io_reg_control_20),
    .io_reg_control_50(qdma_io_reg_control_50),
    .io_reg_control_51(qdma_io_reg_control_51),
    .io_reg_control_52(qdma_io_reg_control_52),
    .io_reg_control_53(qdma_io_reg_control_53),
    .io_reg_control_54(qdma_io_reg_control_54),
    .io_reg_control_55(qdma_io_reg_control_55),
    .io_reg_control_56(qdma_io_reg_control_56),
    .io_reg_control_57(qdma_io_reg_control_57),
    .io_reg_control_58(qdma_io_reg_control_58),
    .io_reg_control_59(qdma_io_reg_control_59),
    .io_reg_control_70(qdma_io_reg_control_70),
    .io_reg_control_71(qdma_io_reg_control_71),
    .io_reg_control_72(qdma_io_reg_control_72),
    .io_reg_control_73(qdma_io_reg_control_73),
    .io_reg_control_74(qdma_io_reg_control_74),
    .io_reg_control_75(qdma_io_reg_control_75),
    .io_reg_control_76(qdma_io_reg_control_76),
    .io_reg_control_77(qdma_io_reg_control_77),
    .io_reg_control_78(qdma_io_reg_control_78),
    .io_reg_control_79(qdma_io_reg_control_79),
    .io_reg_control_80(qdma_io_reg_control_80),
    .io_reg_control_91(qdma_io_reg_control_91),
    .io_reg_control_92(qdma_io_reg_control_92),
    .io_reg_control_93(qdma_io_reg_control_93),
    .io_reg_control_94(qdma_io_reg_control_94),
    .io_reg_status_40(qdma_io_reg_status_40),
    .io_reg_status_51(qdma_io_reg_status_51),
    .io_reg_status_52(qdma_io_reg_status_52),
    .io_reg_status_61(qdma_io_reg_status_61),
    .io_reg_status_71(qdma_io_reg_status_71),
    .io_reg_status_72(qdma_io_reg_status_72),
    .io_reg_status_75(qdma_io_reg_status_75),
    .io_reg_status_76(qdma_io_reg_status_76),
    .io_reg_status_77(qdma_io_reg_status_77),
    .io_reg_status_78(qdma_io_reg_status_78),
    .io_reg_status_79(qdma_io_reg_status_79),
    .io_reg_status_81(qdma_io_reg_status_81),
    .io_axib_aw_ready(qdma_io_axib_aw_ready),
    .io_axib_aw_valid(qdma_io_axib_aw_valid),
    .io_axib_aw_bits_addr(qdma_io_axib_aw_bits_addr),
    .io_axib_aw_bits_burst(qdma_io_axib_aw_bits_burst),
    .io_axib_aw_bits_len(qdma_io_axib_aw_bits_len),
    .io_axib_aw_bits_size(qdma_io_axib_aw_bits_size),
    .io_axib_ar_ready(qdma_io_axib_ar_ready),
    .io_axib_ar_valid(qdma_io_axib_ar_valid),
    .io_axib_ar_bits_addr(qdma_io_axib_ar_bits_addr),
    .io_axib_ar_bits_burst(qdma_io_axib_ar_bits_burst),
    .io_axib_ar_bits_len(qdma_io_axib_ar_bits_len),
    .io_axib_ar_bits_size(qdma_io_axib_ar_bits_size),
    .io_axib_w_ready(qdma_io_axib_w_ready),
    .io_axib_w_valid(qdma_io_axib_w_valid),
    .io_axib_w_bits_data(qdma_io_axib_w_bits_data),
    .io_axib_w_bits_last(qdma_io_axib_w_bits_last),
    .io_axib_w_bits_strb(qdma_io_axib_w_bits_strb),
    .io_axib_r_ready(qdma_io_axib_r_ready),
    .io_axib_r_valid(qdma_io_axib_r_valid),
    .io_axib_r_bits_data(qdma_io_axib_r_bits_data),
    .io_axib_r_bits_last(qdma_io_axib_r_bits_last),
    .io_axib_b_valid(qdma_io_axib_b_valid),
    .io_c2h_status_last(qdma_io_c2h_status_last),
    .io_c2h_status_cmp(qdma_io_c2h_status_cmp),
    .io_c2h_status_valid(qdma_io_c2h_status_valid),
    .io_c2h_status_error(qdma_io_c2h_status_error),
    .io_c2h_status_drop(qdma_io_c2h_status_drop),
    .io_tlb_miss_count(qdma_io_tlb_miss_count)
  );
  h2dcmdqueue h2d_cmd_queue ( // @[Top.scala 86:128]
    .clock(h2d_cmd_queue_clock),
    .reset(h2d_cmd_queue_reset),
    .io_cmd_in_valid(h2d_cmd_queue_io_cmd_in_valid),
    .io_cmd_in_bits_h2c_start_addr(h2d_cmd_queue_io_cmd_in_bits_h2c_start_addr),
    .io_cmd_in_bits_h2m_start_addr(h2d_cmd_queue_io_cmd_in_bits_h2m_start_addr),
    .io_cmd_in_bits_h2m_length(h2d_cmd_queue_io_cmd_in_bits_h2m_length),
    .io_cmd_in_bits_pkt_size(h2d_cmd_queue_io_cmd_in_bits_pkt_size),
    .io_cmd_in_bits_h2c_cpt_addr(h2d_cmd_queue_io_cmd_in_bits_h2c_cpt_addr),
    .io_qin(h2d_cmd_queue_io_qin),
    .io_cmd_out_ready(h2d_cmd_queue_io_cmd_out_ready),
    .io_cmd_out_valid(h2d_cmd_queue_io_cmd_out_valid),
    .io_cmd_out_bits_h2c_start_addr(h2d_cmd_queue_io_cmd_out_bits_h2c_start_addr),
    .io_cmd_out_bits_h2m_start_addr(h2d_cmd_queue_io_cmd_out_bits_h2m_start_addr),
    .io_cmd_out_bits_h2m_length(h2d_cmd_queue_io_cmd_out_bits_h2m_length),
    .io_cmd_out_bits_h2c_cpt_addr(h2d_cmd_queue_io_cmd_out_bits_h2c_cpt_addr),
    .io_h2c_length(h2d_cmd_queue_io_h2c_length),
    .io_h2m_complete(h2d_cmd_queue_io_h2m_complete),
    .io_h2m_cpt_complete(h2d_cmd_queue_io_h2m_cpt_complete),
    .io_last(h2d_cmd_queue_io_last),
    .io_h2m_last(h2d_cmd_queue_io_h2m_last),
    .io_counter(h2d_cmd_queue_io_counter)
  );
  H2C h2c ( // @[Top.scala 98:65]
    .clock(h2c_clock),
    .reset(h2c_reset),
    .io_start_addr(h2c_io_start_addr),
    .io_length(h2c_io_length),
    .io_start(h2c_io_start),
    .io_h2c_cmd_ready(h2c_io_h2c_cmd_ready),
    .io_h2c_cmd_valid(h2c_io_h2c_cmd_valid),
    .io_h2c_cmd_bits_addr(h2c_io_h2c_cmd_bits_addr),
    .io_h2c_cmd_bits_len(h2c_io_h2c_cmd_bits_len),
    .io_complete(h2c_io_complete),
    .io_count_time(h2c_io_count_time),
    .io_send_cmd_count(h2c_io_send_cmd_count)
  );
  d2hcmdqueue d2h_cmd_queue ( // @[Top.scala 111:128]
    .clock(d2h_cmd_queue_clock),
    .reset(d2h_cmd_queue_reset),
    .io_cmd_in_valid(d2h_cmd_queue_io_cmd_in_valid),
    .io_cmd_in_bits_c2h_start_addr(d2h_cmd_queue_io_cmd_in_bits_c2h_start_addr),
    .io_cmd_in_bits_m2h_start_addr(d2h_cmd_queue_io_cmd_in_bits_m2h_start_addr),
    .io_cmd_in_bits_m2h_length(d2h_cmd_queue_io_cmd_in_bits_m2h_length),
    .io_cmd_in_bits_c2h_cpt_addr(d2h_cmd_queue_io_cmd_in_bits_c2h_cpt_addr),
    .io_cmd_in_bits_pkt_size(d2h_cmd_queue_io_cmd_in_bits_pkt_size),
    .io_qin(d2h_cmd_queue_io_qin),
    .io_cmd_out_ready(d2h_cmd_queue_io_cmd_out_ready),
    .io_cmd_out_valid(d2h_cmd_queue_io_cmd_out_valid),
    .io_cmd_out_bits_c2h_start_addr(d2h_cmd_queue_io_cmd_out_bits_c2h_start_addr),
    .io_cmd_out_bits_m2h_start_addr(d2h_cmd_queue_io_cmd_out_bits_m2h_start_addr),
    .io_cmd_out_bits_m2h_length(d2h_cmd_queue_io_cmd_out_bits_m2h_length),
    .io_cmd_out_bits_c2h_cpt_addr(d2h_cmd_queue_io_cmd_out_bits_c2h_cpt_addr),
    .io_c2h_length(d2h_cmd_queue_io_c2h_length),
    .io_m2h_complete(d2h_cmd_queue_io_m2h_complete),
    .io_c2h_finish(d2h_cmd_queue_io_c2h_finish),
    .io_m2h_finish(d2h_cmd_queue_io_m2h_finish),
    .io_m2h_cpt_complete(d2h_cmd_queue_io_m2h_cpt_complete),
    .io_read_count_equal(d2h_cmd_queue_io_read_count_equal),
    .io_empty(d2h_cmd_queue_io_empty),
    .io_h2m_complete_start(d2h_cmd_queue_io_h2m_complete_start),
    .io_h2m_complete(d2h_cmd_queue_io_h2m_complete),
    .io_h2m_cpt_complete(d2h_cmd_queue_io_h2m_cpt_complete),
    .io_m2h_valid_tmpreg(d2h_cmd_queue_io_m2h_valid_tmpreg),
    .io_last(d2h_cmd_queue_io_last),
    .io_counter(d2h_cmd_queue_io_counter)
  );
  C2H c2h ( // @[Top.scala 123:64]
    .clock(c2h_clock),
    .reset(c2h_reset),
    .io_start_addr(c2h_io_start_addr),
    .io_length(c2h_io_length),
    .io_start(c2h_io_start),
    .io_c2h_cmd_ready(c2h_io_c2h_cmd_ready),
    .io_c2h_cmd_valid(c2h_io_c2h_cmd_valid),
    .io_c2h_cmd_bits_addr(c2h_io_c2h_cmd_bits_addr),
    .io_c2h_cmd_bits_pfch_tag(c2h_io_c2h_cmd_bits_pfch_tag),
    .io_c2h_cmd_bits_len(c2h_io_c2h_cmd_bits_len),
    .io_pfch_tag(c2h_io_pfch_tag),
    .io_complete(c2h_io_complete),
    .io_count_time(c2h_io_count_time),
    .io_send_cmd_count(c2h_io_send_cmd_count)
  );
  C2H_Complete c2h_cpt ( // @[Top.scala 137:68]
    .clock(c2h_cpt_clock),
    .reset(c2h_cpt_reset),
    .io_h2c_cpt_addr(c2h_cpt_io_h2c_cpt_addr),
    .io_c2h_cpt_addr(c2h_cpt_io_c2h_cpt_addr),
    .io_p2p_cpt_addr(c2h_cpt_io_p2p_cpt_addr),
    .io_h2c_complete(c2h_cpt_io_h2c_complete),
    .io_c2h_complete(c2h_cpt_io_c2h_complete),
    .io_p2p_complete(c2h_cpt_io_p2p_complete),
    .io_pfch_tag(c2h_cpt_io_pfch_tag),
    .io_h2c_start(c2h_cpt_io_h2c_start),
    .io_c2h_start(c2h_cpt_io_c2h_start),
    .io_h2c_cpt_complete(c2h_cpt_io_h2c_cpt_complete),
    .io_c2h_cpt_complete(c2h_cpt_io_c2h_cpt_complete),
    .io_p2p_cpt_complete(c2h_cpt_io_p2p_cpt_complete),
    .io_polling(c2h_cpt_io_polling),
    .io_c2h_cmd_ready(c2h_cpt_io_c2h_cmd_ready),
    .io_c2h_cmd_valid(c2h_cpt_io_c2h_cmd_valid),
    .io_c2h_cmd_bits_addr(c2h_cpt_io_c2h_cmd_bits_addr),
    .io_c2h_cmd_bits_pfch_tag(c2h_cpt_io_c2h_cmd_bits_pfch_tag),
    .io_c2h_data_ready(c2h_cpt_io_c2h_data_ready),
    .io_c2h_data_valid(c2h_cpt_io_c2h_data_valid)
  );
  H2M h2m ( // @[Top.scala 165:62]
    .clock(h2m_clock),
    .reset(h2m_reset),
    .io_start_addr(h2m_io_start_addr),
    .io_length(h2m_io_length),
    .io_start(h2m_io_start),
    .io_complete(h2m_io_complete),
    .io_awaddr(h2m_io_awaddr),
    .io_awvalid(h2m_io_awvalid),
    .io_awready(h2m_io_awready),
    .io_awlen(h2m_io_awlen),
    .io_wfire(h2m_io_wfire),
    .io_fifo_rden(h2m_io_fifo_rden),
    .io_wlast(h2m_io_wlast),
    .io_last(h2m_io_last),
    .io_clear(h2m_io_clear)
  );
  M2H m2h ( // @[Top.scala 167:62]
    .clock(m2h_clock),
    .reset(m2h_reset),
    .io_start_addr(m2h_io_start_addr),
    .io_length(m2h_io_length),
    .io_start(m2h_io_start),
    .io_complete(m2h_io_complete),
    .io_araddr(m2h_io_araddr),
    .io_arvalid(m2h_io_arvalid),
    .io_arready(m2h_io_arready),
    .io_arlen(m2h_io_arlen),
    .io_rfire(m2h_io_rfire),
    .io_last(m2h_io_last),
    .io_m2h_queue_empty(m2h_io_m2h_queue_empty),
    .io_m2h_valid_tmpreg(m2h_io_m2h_valid_tmpreg),
    .io_read_count_equal(m2h_io_read_count_equal)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(34), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    h2m_start_addr ( // @[CDC.scala 10:25]
    .dest_out(h2m_start_addr_dest_out),
    .dest_clk(h2m_start_addr_dest_clk),
    .src_clk(h2m_start_addr_src_clk),
    .src_in(h2m_start_addr_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(32), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    h2m_length ( // @[CDC.scala 10:25]
    .dest_out(h2m_length_dest_out),
    .dest_clk(h2m_length_dest_clk),
    .src_clk(h2m_length_src_clk),
    .src_in(h2m_length_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4)) h2m_last
     ( // @[CDC.scala 10:25]
    .dest_out(h2m_last_dest_out),
    .dest_clk(h2m_last_dest_clk),
    .src_clk(h2m_last_src_clk),
    .src_in(h2m_last_src_in)
  );
  xpm_cdc_pulse #(.RST_USED(0), .REG_OUTPUT(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4)) h2m_start_pulse
     ( // @[CDC.scala 39:25]
    .dest_pulse(h2m_start_pulse_dest_pulse),
    .dest_clk(h2m_start_pulse_dest_clk),
    .src_clk(h2m_start_pulse_src_clk),
    .src_pulse(h2m_start_pulse_src_pulse)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    h2m_complete ( // @[CDC.scala 10:25]
    .dest_out(h2m_complete_dest_out),
    .dest_clk(h2m_complete_dest_clk),
    .src_clk(h2m_complete_src_clk),
    .src_in(h2m_complete_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4)) h2m_clear
     ( // @[CDC.scala 10:25]
    .dest_out(h2m_clear_dest_out),
    .dest_clk(h2m_clear_dest_clk),
    .src_clk(h2m_clear_src_clk),
    .src_in(h2m_clear_src_in)
  );
  XQueue_34 h2m_cmd_buffer ( // @[XQueue.scala 35:23]
    .clock(h2m_cmd_buffer_clock),
    .reset(h2m_cmd_buffer_reset),
    .io_in_ready(h2m_cmd_buffer_io_in_ready),
    .io_in_valid(h2m_cmd_buffer_io_in_valid),
    .io_in_bits(h2m_cmd_buffer_io_in_bits),
    .io_out_ready(h2m_cmd_buffer_io_out_ready),
    .io_out_valid(h2m_cmd_buffer_io_out_valid),
    .io_out_bits(h2m_cmd_buffer_io_out_bits)
  );
  h2mcmdbufferready h2m_cmd_buffer_ready ( // @[Top.scala 184:120]
    .clock(h2m_cmd_buffer_ready_clock),
    .reset(h2m_cmd_buffer_ready_reset),
    .io_ready(h2m_cmd_buffer_ready_io_ready),
    .io_valid(h2m_cmd_buffer_ready_io_valid),
    .io_complete(h2m_cmd_buffer_ready_io_complete)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(64), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    m2h_start_addr ( // @[CDC.scala 10:25]
    .dest_out(m2h_start_addr_dest_out),
    .dest_clk(m2h_start_addr_dest_clk),
    .src_clk(m2h_start_addr_src_clk),
    .src_in(m2h_start_addr_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(32), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    m2h_length ( // @[CDC.scala 10:25]
    .dest_out(m2h_length_dest_out),
    .dest_clk(m2h_length_dest_clk),
    .src_clk(m2h_length_src_clk),
    .src_in(m2h_length_src_in)
  );
  xpm_cdc_pulse #(.RST_USED(0), .REG_OUTPUT(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4)) m2h_start_pulse
     ( // @[CDC.scala 39:25]
    .dest_pulse(m2h_start_pulse_dest_pulse),
    .dest_clk(m2h_start_pulse_dest_clk),
    .src_clk(m2h_start_pulse_src_clk),
    .src_pulse(m2h_start_pulse_src_pulse)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    m2h_complete ( // @[CDC.scala 10:25]
    .dest_out(m2h_complete_dest_out),
    .dest_clk(m2h_complete_dest_clk),
    .src_clk(m2h_complete_src_clk),
    .src_in(m2h_complete_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4)) m2h_last
     ( // @[CDC.scala 10:25]
    .dest_out(m2h_last_dest_out),
    .dest_clk(m2h_last_dest_clk),
    .src_clk(m2h_last_src_clk),
    .src_in(m2h_last_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    m2h_read_count_equal ( // @[CDC.scala 10:25]
    .dest_out(m2h_read_count_equal_dest_out),
    .dest_clk(m2h_read_count_equal_dest_clk),
    .src_clk(m2h_read_count_equal_src_clk),
    .src_in(m2h_read_count_equal_src_in)
  );
  c2h_status c2h_status ( // @[Top.scala 244:129]
    .clock(c2h_status_clock),
    .reset(c2h_status_reset),
    .io_c2h_start(c2h_status_io_c2h_start),
    .io_c2h_status_last(c2h_status_io_c2h_status_last),
    .io_c2h_status_cmp(c2h_status_io_c2h_status_cmp),
    .io_c2h_status_valid(c2h_status_io_c2h_status_valid),
    .io_c2h_status_error(c2h_status_io_c2h_status_error),
    .io_c2h_status_drop(c2h_status_io_c2h_status_drop),
    .io_c2h_status_last_count(c2h_status_io_c2h_status_last_count),
    .io_c2h_status_cmp_count(c2h_status_io_c2h_status_cmp_count),
    .io_c2h_status_valid_count(c2h_status_io_c2h_status_valid_count),
    .io_c2h_status_error_count(c2h_status_io_c2h_status_error_count),
    .io_c2h_status_drop_count(c2h_status_io_c2h_status_drop_count)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    c2h_status_start ( // @[CDC.scala 10:25]
    .dest_out(c2h_status_start_dest_out),
    .dest_clk(c2h_status_start_dest_clk),
    .src_clk(c2h_status_start_src_clk),
    .src_in(c2h_status_start_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(32), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    last_count ( // @[CDC.scala 10:25]
    .dest_out(last_count_dest_out),
    .dest_clk(last_count_dest_clk),
    .src_clk(last_count_src_clk),
    .src_in(last_count_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(32), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    cmp_count ( // @[CDC.scala 10:25]
    .dest_out(cmp_count_dest_out),
    .dest_clk(cmp_count_dest_clk),
    .src_clk(cmp_count_src_clk),
    .src_in(cmp_count_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(32), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    valid_count ( // @[CDC.scala 10:25]
    .dest_out(valid_count_dest_out),
    .dest_clk(valid_count_dest_clk),
    .src_clk(valid_count_src_clk),
    .src_in(valid_count_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(32), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    error_count ( // @[CDC.scala 10:25]
    .dest_out(error_count_dest_out),
    .dest_clk(error_count_dest_clk),
    .src_clk(error_count_src_clk),
    .src_in(error_count_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(32), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    drop_count ( // @[CDC.scala 10:25]
    .dest_out(drop_count_dest_out),
    .dest_clk(drop_count_dest_clk),
    .src_clk(drop_count_src_clk),
    .src_in(drop_count_src_in)
  );
  xpm_fifo_async
    #(.RD_DATA_COUNT_WIDTH(1), .READ_DATA_WIDTH(256), .USE_ADV_FEATURES("1415"), .WRITE_DATA_WIDTH(512), .FIFO_WRITE_DEPTH(512), .WAKEUP_TIME(0), .PROG_EMPTY_THRESH(10), .READ_MODE("std"), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(1), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("block"), .PROG_FULL_THRESH(10), .FULL_RESET_VALUE(0), .FIFO_READ_LATENCY(1), .DOUT_RESET_VALUE("0"), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    h2m_queue ( // @[Top.scala 275:31]
    .almost_empty(h2m_queue_almost_empty),
    .almost_full(h2m_queue_almost_full),
    .data_valid(h2m_queue_data_valid),
    .dbiterr(h2m_queue_dbiterr),
    .dout(h2m_queue_dout),
    .empty(h2m_queue_empty),
    .full(h2m_queue_full),
    .overflow(h2m_queue_overflow),
    .prog_empty(h2m_queue_prog_empty),
    .prog_full(h2m_queue_prog_full),
    .rd_data_count(h2m_queue_rd_data_count),
    .rd_rst_busy(h2m_queue_rd_rst_busy),
    .sbiterr(h2m_queue_sbiterr),
    .underflow(h2m_queue_underflow),
    .wr_ack(h2m_queue_wr_ack),
    .wr_data_count(h2m_queue_wr_data_count),
    .wr_rst_busy(h2m_queue_wr_rst_busy),
    .din(h2m_queue_din),
    .injectdbiterr(h2m_queue_injectdbiterr),
    .injectsbiterr(h2m_queue_injectsbiterr),
    .rd_clk(h2m_queue_rd_clk),
    .rd_en(h2m_queue_rd_en),
    .rst(h2m_queue_rst),
    .sleep(h2m_queue_sleep),
    .wr_clk(h2m_queue_wr_clk),
    .wr_en(h2m_queue_wr_en)
  );
  xpm_fifo_async
    #(.RD_DATA_COUNT_WIDTH(1), .READ_DATA_WIDTH(512), .USE_ADV_FEATURES("1415"), .WRITE_DATA_WIDTH(256), .FIFO_WRITE_DEPTH(512), .WAKEUP_TIME(0), .PROG_EMPTY_THRESH(10), .READ_MODE("std"), .SIM_ASSERT_CHK(0), .WR_DATA_COUNT_WIDTH(1), .ECC_MODE("no_ecc"), .FIFO_MEMORY_TYPE("block"), .PROG_FULL_THRESH(10), .FULL_RESET_VALUE(0), .FIFO_READ_LATENCY(1), .DOUT_RESET_VALUE("0"), .RELATED_CLOCKS(0), .CASCADE_HEIGHT(0), .CDC_SYNC_STAGES(2))
    m2h_queue_ ( // @[Top.scala 276:31]
    .almost_empty(m2h_queue__almost_empty),
    .almost_full(m2h_queue__almost_full),
    .data_valid(m2h_queue__data_valid),
    .dbiterr(m2h_queue__dbiterr),
    .dout(m2h_queue__dout),
    .empty(m2h_queue__empty),
    .full(m2h_queue__full),
    .overflow(m2h_queue__overflow),
    .prog_empty(m2h_queue__prog_empty),
    .prog_full(m2h_queue__prog_full),
    .rd_data_count(m2h_queue__rd_data_count),
    .rd_rst_busy(m2h_queue__rd_rst_busy),
    .sbiterr(m2h_queue__sbiterr),
    .underflow(m2h_queue__underflow),
    .wr_ack(m2h_queue__wr_ack),
    .wr_data_count(m2h_queue__wr_data_count),
    .wr_rst_busy(m2h_queue__wr_rst_busy),
    .din(m2h_queue__din),
    .injectdbiterr(m2h_queue__injectdbiterr),
    .injectsbiterr(m2h_queue__injectsbiterr),
    .rd_clk(m2h_queue__rd_clk),
    .rd_en(m2h_queue__rd_en),
    .rst(m2h_queue__rst),
    .sleep(m2h_queue__sleep),
    .wr_clk(m2h_queue__wr_clk),
    .wr_en(m2h_queue__wr_en)
  );
  validreg h2m_valid_tmpreg ( // @[Top.scala 289:118]
    .clock(h2m_valid_tmpreg_clock),
    .reset(h2m_valid_tmpreg_reset),
    .io_ready(h2m_valid_tmpreg_io_ready),
    .io_valid(h2m_valid_tmpreg_io_valid),
    .io_tmpreg(h2m_valid_tmpreg_io_tmpreg)
  );
  validreg m2h_valid_tmpreg ( // @[Top.scala 305:120]
    .clock(m2h_valid_tmpreg_clock),
    .reset(m2h_valid_tmpreg_reset),
    .io_ready(m2h_valid_tmpreg_io_ready),
    .io_valid(m2h_valid_tmpreg_io_valid),
    .io_tmpreg(m2h_valid_tmpreg_io_tmpreg)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    m2h_queue_empty ( // @[CDC.scala 10:25]
    .dest_out(m2h_queue_empty_dest_out),
    .dest_clk(m2h_queue_empty_dest_clk),
    .src_clk(m2h_queue_empty_src_clk),
    .src_in(m2h_queue_empty_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    m2h_valid_tmpreg_tom2h ( // @[CDC.scala 10:25]
    .dest_out(m2h_valid_tmpreg_tom2h_dest_out),
    .dest_clk(m2h_valid_tmpreg_tom2h_dest_clk),
    .src_clk(m2h_valid_tmpreg_tom2h_src_clk),
    .src_in(m2h_valid_tmpreg_tom2h_src_in)
  );
  AXIClockConverterBlackBox axicc ( // @[Top.scala 356:27]
    .s_axi_awaddr(axicc_s_axi_awaddr),
    .s_axi_awlen(axicc_s_axi_awlen),
    .s_axi_awsize(axicc_s_axi_awsize),
    .s_axi_awburst(axicc_s_axi_awburst),
    .s_axi_awlock(axicc_s_axi_awlock),
    .s_axi_awcache(axicc_s_axi_awcache),
    .s_axi_awprot(axicc_s_axi_awprot),
    .s_axi_awregion(axicc_s_axi_awregion),
    .s_axi_awqos(axicc_s_axi_awqos),
    .s_axi_awvalid(axicc_s_axi_awvalid),
    .s_axi_awready(axicc_s_axi_awready),
    .s_axi_wdata(axicc_s_axi_wdata),
    .s_axi_wstrb(axicc_s_axi_wstrb),
    .s_axi_wlast(axicc_s_axi_wlast),
    .s_axi_wvalid(axicc_s_axi_wvalid),
    .s_axi_wready(axicc_s_axi_wready),
    .s_axi_bresp(axicc_s_axi_bresp),
    .s_axi_bvalid(axicc_s_axi_bvalid),
    .s_axi_bready(axicc_s_axi_bready),
    .s_axi_araddr(axicc_s_axi_araddr),
    .s_axi_arlen(axicc_s_axi_arlen),
    .s_axi_arsize(axicc_s_axi_arsize),
    .s_axi_arburst(axicc_s_axi_arburst),
    .s_axi_arlock(axicc_s_axi_arlock),
    .s_axi_arcache(axicc_s_axi_arcache),
    .s_axi_arprot(axicc_s_axi_arprot),
    .s_axi_arregion(axicc_s_axi_arregion),
    .s_axi_arqos(axicc_s_axi_arqos),
    .s_axi_arvalid(axicc_s_axi_arvalid),
    .s_axi_arready(axicc_s_axi_arready),
    .s_axi_rdata(axicc_s_axi_rdata),
    .s_axi_rresp(axicc_s_axi_rresp),
    .s_axi_rlast(axicc_s_axi_rlast),
    .s_axi_rvalid(axicc_s_axi_rvalid),
    .s_axi_rready(axicc_s_axi_rready),
    .s_axi_aclk(axicc_s_axi_aclk),
    .s_axi_aresetn(axicc_s_axi_aresetn),
    .m_axi_aclk(axicc_m_axi_aclk),
    .m_axi_aresetn(axicc_m_axi_aresetn),
    .m_axi_awaddr(axicc_m_axi_awaddr),
    .m_axi_awlen(axicc_m_axi_awlen),
    .m_axi_awsize(axicc_m_axi_awsize),
    .m_axi_awburst(axicc_m_axi_awburst),
    .m_axi_awlock(axicc_m_axi_awlock),
    .m_axi_awcache(axicc_m_axi_awcache),
    .m_axi_awprot(axicc_m_axi_awprot),
    .m_axi_awregion(axicc_m_axi_awregion),
    .m_axi_awqos(axicc_m_axi_awqos),
    .m_axi_awvalid(axicc_m_axi_awvalid),
    .m_axi_awready(axicc_m_axi_awready),
    .m_axi_wdata(axicc_m_axi_wdata),
    .m_axi_wstrb(axicc_m_axi_wstrb),
    .m_axi_wlast(axicc_m_axi_wlast),
    .m_axi_wvalid(axicc_m_axi_wvalid),
    .m_axi_wready(axicc_m_axi_wready),
    .m_axi_bresp(axicc_m_axi_bresp),
    .m_axi_bvalid(axicc_m_axi_bvalid),
    .m_axi_bready(axicc_m_axi_bready),
    .m_axi_araddr(axicc_m_axi_araddr),
    .m_axi_arlen(axicc_m_axi_arlen),
    .m_axi_arsize(axicc_m_axi_arsize),
    .m_axi_arburst(axicc_m_axi_arburst),
    .m_axi_arlock(axicc_m_axi_arlock),
    .m_axi_arcache(axicc_m_axi_arcache),
    .m_axi_arprot(axicc_m_axi_arprot),
    .m_axi_arregion(axicc_m_axi_arregion),
    .m_axi_arqos(axicc_m_axi_arqos),
    .m_axi_arvalid(axicc_m_axi_arvalid),
    .m_axi_arready(axicc_m_axi_arready),
    .m_axi_rdata(axicc_m_axi_rdata),
    .m_axi_rresp(axicc_m_axi_rresp),
    .m_axi_rlast(axicc_m_axi_rlast),
    .m_axi_rvalid(axicc_m_axi_rvalid),
    .m_axi_rready(axicc_m_axi_rready)
  );
  AXIDataWidthConverterBlackBox axidwc ( // @[Top.scala 404:28]
    .s_axi_awaddr(axidwc_s_axi_awaddr),
    .s_axi_awlen(axidwc_s_axi_awlen),
    .s_axi_awsize(axidwc_s_axi_awsize),
    .s_axi_awburst(axidwc_s_axi_awburst),
    .s_axi_awlock(axidwc_s_axi_awlock),
    .s_axi_awcache(axidwc_s_axi_awcache),
    .s_axi_awprot(axidwc_s_axi_awprot),
    .s_axi_awregion(axidwc_s_axi_awregion),
    .s_axi_awqos(axidwc_s_axi_awqos),
    .s_axi_awvalid(axidwc_s_axi_awvalid),
    .s_axi_awready(axidwc_s_axi_awready),
    .s_axi_wdata(axidwc_s_axi_wdata),
    .s_axi_wstrb(axidwc_s_axi_wstrb),
    .s_axi_wlast(axidwc_s_axi_wlast),
    .s_axi_wvalid(axidwc_s_axi_wvalid),
    .s_axi_wready(axidwc_s_axi_wready),
    .s_axi_bresp(axidwc_s_axi_bresp),
    .s_axi_bvalid(axidwc_s_axi_bvalid),
    .s_axi_bready(axidwc_s_axi_bready),
    .s_axi_araddr(axidwc_s_axi_araddr),
    .s_axi_arlen(axidwc_s_axi_arlen),
    .s_axi_arsize(axidwc_s_axi_arsize),
    .s_axi_arburst(axidwc_s_axi_arburst),
    .s_axi_arlock(axidwc_s_axi_arlock),
    .s_axi_arcache(axidwc_s_axi_arcache),
    .s_axi_arprot(axidwc_s_axi_arprot),
    .s_axi_arregion(axidwc_s_axi_arregion),
    .s_axi_arqos(axidwc_s_axi_arqos),
    .s_axi_arvalid(axidwc_s_axi_arvalid),
    .s_axi_arready(axidwc_s_axi_arready),
    .s_axi_rdata(axidwc_s_axi_rdata),
    .s_axi_rresp(axidwc_s_axi_rresp),
    .s_axi_rlast(axidwc_s_axi_rlast),
    .s_axi_rvalid(axidwc_s_axi_rvalid),
    .s_axi_rready(axidwc_s_axi_rready),
    .s_axi_aclk(axidwc_s_axi_aclk),
    .s_axi_aresetn(axidwc_s_axi_aresetn),
    .m_axi_awaddr(axidwc_m_axi_awaddr),
    .m_axi_awlen(axidwc_m_axi_awlen),
    .m_axi_awsize(axidwc_m_axi_awsize),
    .m_axi_awburst(axidwc_m_axi_awburst),
    .m_axi_awlock(axidwc_m_axi_awlock),
    .m_axi_awcache(axidwc_m_axi_awcache),
    .m_axi_awprot(axidwc_m_axi_awprot),
    .m_axi_awregion(axidwc_m_axi_awregion),
    .m_axi_awqos(axidwc_m_axi_awqos),
    .m_axi_awvalid(axidwc_m_axi_awvalid),
    .m_axi_awready(axidwc_m_axi_awready),
    .m_axi_wdata(axidwc_m_axi_wdata),
    .m_axi_wstrb(axidwc_m_axi_wstrb),
    .m_axi_wlast(axidwc_m_axi_wlast),
    .m_axi_wvalid(axidwc_m_axi_wvalid),
    .m_axi_wready(axidwc_m_axi_wready),
    .m_axi_bresp(axidwc_m_axi_bresp),
    .m_axi_bvalid(axidwc_m_axi_bvalid),
    .m_axi_bready(axidwc_m_axi_bready),
    .m_axi_araddr(axidwc_m_axi_araddr),
    .m_axi_arlen(axidwc_m_axi_arlen),
    .m_axi_arsize(axidwc_m_axi_arsize),
    .m_axi_arburst(axidwc_m_axi_arburst),
    .m_axi_arlock(axidwc_m_axi_arlock),
    .m_axi_arcache(axidwc_m_axi_arcache),
    .m_axi_arprot(axidwc_m_axi_arprot),
    .m_axi_arregion(axidwc_m_axi_arregion),
    .m_axi_arqos(axidwc_m_axi_arqos),
    .m_axi_arvalid(axidwc_m_axi_arvalid),
    .m_axi_arready(axidwc_m_axi_arready),
    .m_axi_rdata(axidwc_m_axi_rdata),
    .m_axi_rresp(axidwc_m_axi_rresp),
    .m_axi_rlast(axidwc_m_axi_rlast),
    .m_axi_rvalid(axidwc_m_axi_rvalid),
    .m_axi_rready(axidwc_m_axi_rready)
  );
  p2p_counter p2p_counter ( // @[Top.scala 472:102]
    .clock(p2p_counter_clock),
    .reset(p2p_counter_reset),
    .io_start(p2p_counter_io_start),
    .io_length(p2p_counter_io_length),
    .io_wready(p2p_counter_io_wready),
    .io_wvalid(p2p_counter_io_wvalid),
    .io_wdatasample(p2p_counter_io_wdatasample),
    .io_p2p_complete(p2p_counter_io_p2p_complete),
    .io_p2p_cpt_complete(p2p_counter_io_p2p_cpt_complete)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(64), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    p2p_cpt_addr ( // @[CDC.scala 10:25]
    .dest_out(p2p_cpt_addr_dest_out),
    .dest_clk(p2p_cpt_addr_dest_clk),
    .src_clk(p2p_cpt_addr_src_clk),
    .src_in(p2p_cpt_addr_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(32), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4))
    p2p_length ( // @[CDC.scala 10:25]
    .dest_out(p2p_length_dest_out),
    .dest_clk(p2p_length_dest_clk),
    .src_clk(p2p_length_src_clk),
    .src_in(p2p_length_src_in)
  );
  xpm_cdc_array_single #(.SRC_INPUT_REG(1), .WIDTH(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4)) p2p_start
     ( // @[CDC.scala 10:25]
    .dest_out(p2p_start_dest_out),
    .dest_clk(p2p_start_dest_clk),
    .src_clk(p2p_start_src_clk),
    .src_in(p2p_start_src_in)
  );
  xpm_cdc_pulse #(.RST_USED(0), .REG_OUTPUT(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4)) p2p_complete ( // @[CDC.scala 39:25]
    .dest_pulse(p2p_complete_dest_pulse),
    .dest_clk(p2p_complete_dest_clk),
    .src_clk(p2p_complete_src_clk),
    .src_pulse(p2p_complete_src_pulse)
  );
  xpm_cdc_pulse #(.RST_USED(0), .REG_OUTPUT(1), .SIM_ASSERT_CHK(0), .INIT_SYNC_FF(0), .DEST_SYNC_FF(4)) p2p_cpt_complete
     ( // @[CDC.scala 39:25]
    .dest_pulse(p2p_cpt_complete_dest_pulse),
    .dest_clk(p2p_cpt_complete_dest_clk),
    .src_clk(p2p_cpt_complete_src_clk),
    .src_pulse(p2p_cpt_complete_src_pulse)
  );
  assign qdma_pin_tx_p = qdma_io_pin_tx_p; // @[Top.scala 58:21]
  assign qdma_pin_tx_n = qdma_io_pin_tx_n; // @[Top.scala 58:21]
  assign mmcm_io_CLKIN1 = mmcm_io_CLKIN1_pad_O; // @[Top.scala 26:25]
  assign mmcm_io_CLKIN1_pad_I = sys_100M_0_p; // @[Buf.scala 52:26]
  assign mmcm_io_CLKIN1_pad_IB = sys_100M_0_n; // @[Buf.scala 53:27]
  assign hbmDriver_clock = mmcm_io_CLKOUT0;
  assign hbmDriver_io_axi_hbm_0_aw_valid = h2m_io_awvalid; // @[Top.scala 328:81]
  assign hbmDriver_io_axi_hbm_0_aw_bits_addr = h2m_io_awaddr; // @[Top.scala 327:81]
  assign hbmDriver_io_axi_hbm_0_aw_bits_len = h2m_io_awlen[3:0]; // @[Top.scala 331:81]
  assign hbmDriver_io_axi_hbm_0_ar_valid = m2h_io_arvalid; // @[Top.scala 343:81]
  assign hbmDriver_io_axi_hbm_0_ar_bits_addr = m2h_io_araddr; // @[Top.scala 342:81]
  assign hbmDriver_io_axi_hbm_0_ar_bits_len = m2h_io_arlen[3:0]; // @[Top.scala 347:81]
  assign hbmDriver_io_axi_hbm_0_w_valid = h2m_io_fifo_rden & h2m_queue_data_valid + h2m_valid_tmpreg_io_tmpreg; // @[Top.scala 292:71]
  assign hbmDriver_io_axi_hbm_0_w_bits_data = h2m_queue_dout; // @[Top.scala 288:81]
  assign hbmDriver_io_axi_hbm_0_w_bits_last = h2m_io_wlast; // @[Top.scala 323:81]
  assign hbmDriver_io_axi_hbm_0_r_ready = ~m2h_queue__almost_full & ~m2h_queue__full; // @[Top.scala 300:94]
  assign hbmDriver_io_axi_hbm_1_aw_valid = axidwc_m_axi_awvalid; // @[Top.scala 451:41]
  assign hbmDriver_io_axi_hbm_1_aw_bits_addr = axidwc_m_axi_awaddr; // @[Top.scala 447:41]
  assign hbmDriver_io_axi_hbm_1_aw_bits_burst = axidwc_m_axi_awburst; // @[Top.scala 450:41]
  assign hbmDriver_io_axi_hbm_1_aw_bits_len = axidwc_m_axi_awlen[3:0]; // @[Top.scala 448:41]
  assign hbmDriver_io_axi_hbm_1_aw_bits_size = axidwc_m_axi_awsize; // @[Top.scala 449:41]
  assign hbmDriver_io_axi_hbm_1_ar_valid = axidwc_m_axi_arvalid; // @[Top.scala 462:41]
  assign hbmDriver_io_axi_hbm_1_ar_bits_addr = axidwc_m_axi_araddr; // @[Top.scala 458:41]
  assign hbmDriver_io_axi_hbm_1_ar_bits_burst = axidwc_m_axi_arburst; // @[Top.scala 461:41]
  assign hbmDriver_io_axi_hbm_1_ar_bits_len = axidwc_m_axi_arlen[3:0]; // @[Top.scala 459:41]
  assign hbmDriver_io_axi_hbm_1_ar_bits_size = axidwc_m_axi_arsize; // @[Top.scala 460:41]
  assign hbmDriver_io_axi_hbm_1_w_valid = axidwc_m_axi_wvalid; // @[Top.scala 456:41]
  assign hbmDriver_io_axi_hbm_1_w_bits_data = axidwc_m_axi_wdata; // @[Top.scala 453:41]
  assign hbmDriver_io_axi_hbm_1_w_bits_last = axidwc_m_axi_wlast; // @[Top.scala 455:41]
  assign hbmDriver_io_axi_hbm_1_w_bits_strb = axidwc_m_axi_wstrb; // @[Top.scala 454:41]
  assign hbmDriver_io_axi_hbm_1_r_ready = axidwc_m_axi_rready; // @[Top.scala 467:41]
  assign hbmDriver_io_axi_hbm_1_b_ready = axidwc_m_axi_bready; // @[Top.scala 469:49]
  assign qdma_io_pin_rx_p = qdma_pin_rx_p; // @[Top.scala 58:21]
  assign qdma_io_pin_rx_n = qdma_pin_rx_n; // @[Top.scala 58:21]
  assign qdma_io_pin_sys_clk_p = qdma_pin_sys_clk_p; // @[Top.scala 58:21]
  assign qdma_io_pin_sys_clk_n = qdma_pin_sys_clk_n; // @[Top.scala 58:21]
  assign qdma_io_pin_sys_rst_n = qdma_pin_sys_rst_n; // @[Top.scala 58:21]
  assign qdma_io_user_clk = mmcm_io_CLKOUT1; // @[Top.scala 60:33]
  assign qdma_io_user_arstn = mmcm_io_LOCKED; // @[Top.scala 61:33]
  assign qdma_io_h2c_cmd_valid = h2c_io_h2c_cmd_valid; // @[Top.scala 103:81]
  assign qdma_io_h2c_cmd_bits_addr = h2c_io_h2c_cmd_bits_addr; // @[Top.scala 103:81]
  assign qdma_io_h2c_cmd_bits_len = h2c_io_h2c_cmd_bits_len; // @[Top.scala 103:81]
  assign qdma_io_h2c_data_ready = ~h2m_queue_almost_full & ~h2m_queue_full; // @[Top.scala 284:102]
  assign qdma_io_c2h_cmd_valid = c2h_cpt_io_c2h_cmd_valid ? c2h_cpt_io_c2h_cmd_valid : c2h_io_c2h_cmd_valid; // @[Top.scala 155:79]
  assign qdma_io_c2h_cmd_bits_addr = c2h_cpt_io_c2h_cmd_valid ? c2h_cpt_io_c2h_cmd_bits_addr : c2h_io_c2h_cmd_bits_addr; // @[Top.scala 156:79]
  assign qdma_io_c2h_cmd_bits_pfch_tag = c2h_cpt_io_c2h_cmd_valid ? c2h_cpt_io_c2h_cmd_bits_pfch_tag :
    c2h_io_c2h_cmd_bits_pfch_tag; // @[Top.scala 156:79]
  assign qdma_io_c2h_cmd_bits_len = c2h_cpt_io_c2h_cmd_valid ? 32'h40 : c2h_io_c2h_cmd_bits_len; // @[Top.scala 156:79]
  assign qdma_io_c2h_data_valid = c2h_cpt_io_c2h_data_valid ? c2h_cpt_io_c2h_data_valid : m2h_queue__data_valid +
    m2h_valid_tmpreg_io_tmpreg; // @[Top.scala 308:79]
  assign qdma_io_c2h_data_bits_data = c2h_cpt_io_c2h_data_valid ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff
     : m2h_queue__dout; // @[Top.scala 304:79]
  assign qdma_io_reg_status_40 = qdma_io_tlb_miss_count; // @[Top.scala 268:73]
  assign qdma_io_reg_status_51 = h2c_io_count_time; // @[Top.scala 105:81]
  assign qdma_io_reg_status_52 = h2c_io_send_cmd_count; // @[Top.scala 106:73]
  assign qdma_io_reg_status_61 = h2d_cmd_queue_io_counter; // @[Top.scala 239:34]
  assign qdma_io_reg_status_71 = c2h_io_count_time; // @[Top.scala 131:81]
  assign qdma_io_reg_status_72 = c2h_io_send_cmd_count; // @[Top.scala 132:73]
  assign qdma_io_reg_status_75 = last_count_dest_out; // @[Top.scala 259:73]
  assign qdma_io_reg_status_76 = cmp_count_dest_out; // @[Top.scala 261:73]
  assign qdma_io_reg_status_77 = valid_count_dest_out; // @[Top.scala 263:73]
  assign qdma_io_reg_status_78 = error_count_dest_out; // @[Top.scala 265:73]
  assign qdma_io_reg_status_79 = drop_count_dest_out; // @[Top.scala 267:73]
  assign qdma_io_reg_status_81 = d2h_cmd_queue_io_counter; // @[Top.scala 240:34]
  assign qdma_io_axib_aw_ready = axicc_s_axi_awready; // @[Top.scala 367:57]
  assign qdma_io_axib_ar_ready = axicc_s_axi_arready; // @[Top.scala 378:57]
  assign qdma_io_axib_w_ready = axicc_s_axi_wready; // @[Top.scala 372:57]
  assign qdma_io_axib_r_valid = axicc_s_axi_rvalid; // @[Top.scala 381:57]
  assign qdma_io_axib_r_bits_data = axicc_s_axi_rdata; // @[Top.scala 379:57]
  assign qdma_io_axib_r_bits_last = axicc_s_axi_rlast; // @[Top.scala 380:57]
  assign qdma_io_axib_b_valid = axicc_s_axi_bvalid; // @[Top.scala 383:57]
  assign h2d_cmd_queue_clock = mmcm_io_CLKOUT1;
  assign h2d_cmd_queue_reset = ~mmcm_io_LOCKED; // @[Top.scala 86:110]
  assign h2d_cmd_queue_io_cmd_in_valid = h2d_cmd_queue_io_cmd_in_valid_REG_2 & ~h2d_cmd_queue_io_cmd_in_valid_REG_3; // @[Top.scala 37:37]
  assign h2d_cmd_queue_io_cmd_in_bits_h2c_start_addr = {qdma_io_reg_control_50,qdma_io_reg_control_51}; // @[Cat.scala 30:58]
  assign h2d_cmd_queue_io_cmd_in_bits_h2m_start_addr = {qdma_io_reg_control_52[1:0],qdma_io_reg_control_53}; // @[Cat.scala 30:58]
  assign h2d_cmd_queue_io_cmd_in_bits_h2m_length = qdma_io_reg_control_54; // @[Top.scala 91:57]
  assign h2d_cmd_queue_io_cmd_in_bits_pkt_size = qdma_io_reg_control_55; // @[Top.scala 92:57]
  assign h2d_cmd_queue_io_cmd_in_bits_h2c_cpt_addr = {qdma_io_reg_control_57,qdma_io_reg_control_58}; // @[Cat.scala 30:58]
  assign h2d_cmd_queue_io_qin = qdma_io_reg_control_56; // @[Top.scala 93:73]
  assign h2d_cmd_queue_io_cmd_out_ready = h2c_io_complete & h2m_cmd_buffer_io_in_ready & (~h2d_cmd_queue_io_last |
    h2d_cmd_queue_io_last & h2m_clear_dest_out); // @[Top.scala 209:113]
  assign h2d_cmd_queue_io_h2m_cpt_complete = c2h_cpt_io_h2c_cpt_complete; // @[Top.scala 145:73]
  assign h2c_clock = mmcm_io_CLKOUT1;
  assign h2c_reset = ~mmcm_io_LOCKED; // @[Top.scala 98:47]
  assign h2c_io_start_addr = h2d_cmd_queue_io_cmd_out_bits_h2c_start_addr; // @[Top.scala 100:81]
  assign h2c_io_length = h2d_cmd_queue_io_h2c_length; // @[Top.scala 101:81]
  assign h2c_io_start = h2d_cmd_queue_io_cmd_out_ready & h2d_cmd_queue_io_cmd_out_valid; // @[Decoupled.scala 40:37]
  assign h2c_io_h2c_cmd_ready = qdma_io_h2c_cmd_ready; // @[Top.scala 103:81]
  assign d2h_cmd_queue_clock = mmcm_io_CLKOUT1;
  assign d2h_cmd_queue_reset = ~mmcm_io_LOCKED; // @[Top.scala 111:110]
  assign d2h_cmd_queue_io_cmd_in_valid = d2h_cmd_queue_io_cmd_in_valid_REG_2 & ~d2h_cmd_queue_io_cmd_in_valid_REG_3; // @[Top.scala 37:37]
  assign d2h_cmd_queue_io_cmd_in_bits_c2h_start_addr = {qdma_io_reg_control_70,qdma_io_reg_control_71}; // @[Cat.scala 30:58]
  assign d2h_cmd_queue_io_cmd_in_bits_m2h_start_addr = {qdma_io_reg_control_72[1:0],qdma_io_reg_control_73}; // @[Cat.scala 30:58]
  assign d2h_cmd_queue_io_cmd_in_bits_m2h_length = qdma_io_reg_control_74; // @[Top.scala 116:57]
  assign d2h_cmd_queue_io_cmd_in_bits_c2h_cpt_addr = {qdma_io_reg_control_77,qdma_io_reg_control_78}; // @[Cat.scala 30:58]
  assign d2h_cmd_queue_io_cmd_in_bits_pkt_size = qdma_io_reg_control_75; // @[Top.scala 117:57]
  assign d2h_cmd_queue_io_qin = qdma_io_reg_control_76; // @[Top.scala 118:73]
  assign d2h_cmd_queue_io_cmd_out_ready = c2h_io_complete & m2h_complete_dest_out & c2h_cpt_io_c2h_cpt_complete; // @[Top.scala 227:111]
  assign d2h_cmd_queue_io_c2h_finish = c2h_io_complete; // @[Top.scala 228:73]
  assign d2h_cmd_queue_io_m2h_finish = m2h_complete_dest_out; // @[Top.scala 229:73]
  assign d2h_cmd_queue_io_m2h_cpt_complete = c2h_cpt_io_c2h_cpt_complete; // @[Top.scala 150:73]
  assign d2h_cmd_queue_io_read_count_equal = m2h_read_count_equal_dest_out; // @[Top.scala 237:65]
  assign d2h_cmd_queue_io_empty = m2h_queue__empty; // @[Top.scala 310:73]
  assign d2h_cmd_queue_io_h2m_complete_start = h2d_cmd_queue_io_h2m_complete & ~d2h_cmd_queue_io_h2m_complete_start_REG; // @[Top.scala 37:37]
  assign d2h_cmd_queue_io_h2m_cpt_complete = c2h_cpt_io_h2c_cpt_complete; // @[Top.scala 146:73]
  assign d2h_cmd_queue_io_m2h_valid_tmpreg = m2h_valid_tmpreg_io_tmpreg; // @[Top.scala 317:65]
  assign c2h_clock = mmcm_io_CLKOUT1;
  assign c2h_reset = ~mmcm_io_LOCKED; // @[Top.scala 123:46]
  assign c2h_io_start_addr = d2h_cmd_queue_io_cmd_out_bits_c2h_start_addr; // @[Top.scala 126:81]
  assign c2h_io_length = d2h_cmd_queue_io_c2h_length; // @[Top.scala 127:81]
  assign c2h_io_start = d2h_cmd_queue_io_cmd_out_ready & d2h_cmd_queue_io_cmd_out_valid; // @[Decoupled.scala 40:37]
  assign c2h_io_c2h_cmd_ready = qdma_io_c2h_cmd_ready & ~c2h_cpt_io_c2h_cmd_valid; // @[Top.scala 157:98]
  assign c2h_io_pfch_tag = qdma_io_reg_control_80; // @[Top.scala 129:81]
  assign c2h_cpt_clock = mmcm_io_CLKOUT1;
  assign c2h_cpt_reset = ~mmcm_io_LOCKED; // @[Top.scala 137:50]
  assign c2h_cpt_io_h2c_cpt_addr = h2d_cmd_queue_io_cmd_out_bits_h2c_cpt_addr; // @[Top.scala 144:73]
  assign c2h_cpt_io_c2h_cpt_addr = d2h_cmd_queue_io_cmd_out_bits_c2h_cpt_addr; // @[Top.scala 149:73]
  assign c2h_cpt_io_p2p_cpt_addr = {qdma_io_reg_control_92,qdma_io_reg_control_93}; // @[Cat.scala 30:58]
  assign c2h_cpt_io_h2c_complete = d2h_cmd_queue_io_h2m_complete; // @[Top.scala 143:73]
  assign c2h_cpt_io_c2h_complete = d2h_cmd_queue_io_m2h_complete; // @[Top.scala 148:73]
  assign c2h_cpt_io_p2p_complete = p2p_complete_dest_pulse; // @[Top.scala 492:49]
  assign c2h_cpt_io_pfch_tag = qdma_io_reg_control_80; // @[Top.scala 151:81]
  assign c2h_cpt_io_h2c_start = h2d_cmd_queue_io_last & ~c2h_cpt_io_h2c_start_REG; // @[Top.scala 37:37]
  assign c2h_cpt_io_c2h_start = d2h_cmd_queue_io_last & ~c2h_cpt_io_c2h_start_REG; // @[Top.scala 37:37]
  assign c2h_cpt_io_polling = qdma_io_reg_control_20; // @[Top.scala 140:81]
  assign c2h_cpt_io_c2h_cmd_ready = qdma_io_c2h_cmd_ready; // @[Top.scala 158:73]
  assign c2h_cpt_io_c2h_data_ready = qdma_io_c2h_data_ready; // @[Top.scala 159:73]
  assign h2m_clock = hbmDriver_io_hbm_clk;
  assign h2m_reset = ~hbm_rstn; // @[Top.scala 165:45]
  assign h2m_io_start_addr = h2m_start_addr_dest_out; // @[Top.scala 201:73]
  assign h2m_io_length = h2m_length_dest_out; // @[Top.scala 202:73]
  assign h2m_io_start = h2m_io_start_REG; // @[Top.scala 206:81]
  assign h2m_io_awready = hbmDriver_io_axi_hbm_0_aw_ready; // @[Top.scala 329:81]
  assign h2m_io_wfire = hbmDriver_io_axi_hbm_0_w_ready & hbmDriver_io_axi_hbm_0_w_valid; // @[Decoupled.scala 40:37]
  assign h2m_io_last = h2m_last_dest_out; // @[Top.scala 203:73]
  assign m2h_clock = hbmDriver_io_hbm_clk;
  assign m2h_reset = ~hbm_rstn; // @[Top.scala 167:45]
  assign m2h_io_start_addr = m2h_start_addr_dest_out[33:0]; // @[Top.scala 222:73]
  assign m2h_io_length = m2h_length_dest_out; // @[Top.scala 223:73]
  assign m2h_io_start = m2h_io_start_REG; // @[Top.scala 224:81]
  assign m2h_io_arready = hbmDriver_io_axi_hbm_0_ar_ready; // @[Top.scala 344:81]
  assign m2h_io_rfire = hbmDriver_io_axi_hbm_0_r_ready & hbmDriver_io_axi_hbm_0_r_valid; // @[Decoupled.scala 40:37]
  assign m2h_io_last = m2h_last_dest_out; // @[Top.scala 234:73]
  assign m2h_io_m2h_queue_empty = m2h_queue_empty_dest_out; // @[Top.scala 313:73]
  assign m2h_io_m2h_valid_tmpreg = m2h_valid_tmpreg_tom2h_dest_out; // @[Top.scala 316:73]
  assign h2m_start_addr_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign h2m_start_addr_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign h2m_start_addr_src_in = h2m_start_addr_reg; // @[Top.scala 197:73]
  assign h2m_length_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign h2m_length_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign h2m_length_src_in = h2m_length_reg[31:0]; // @[Top.scala 198:73]
  assign h2m_last_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign h2m_last_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign h2m_last_src_in = h2m_last_reg; // @[Top.scala 199:81]
  assign h2m_start_pulse_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 41:29]
  assign h2m_start_pulse_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 40:29]
  assign h2m_start_pulse_src_pulse = h2m_cmd_buffer_io_out_ready & h2m_cmd_buffer_io_out_valid; // @[Decoupled.scala 40:37]
  assign h2m_complete_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign h2m_complete_src_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 11:28]
  assign h2m_complete_src_in = h2m_io_complete; // @[Top.scala 176:73]
  assign h2m_clear_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign h2m_clear_src_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 11:28]
  assign h2m_clear_src_in = h2m_io_clear; // @[Top.scala 178:81]
  assign h2m_cmd_buffer_clock = mmcm_io_CLKOUT1;
  assign h2m_cmd_buffer_reset = ~mmcm_io_LOCKED; // @[Top.scala 180:110]
  assign h2m_cmd_buffer_io_in_valid = h2d_cmd_queue_io_cmd_out_ready & h2d_cmd_queue_io_cmd_out_valid; // @[Decoupled.scala 40:37]
  assign h2m_cmd_buffer_io_in_bits = {h2m_cmd_buffer_io_in_bits_hi,h2d_cmd_queue_io_cmd_out_bits_h2m_length}; // @[Cat.scala 30:58]
  assign h2m_cmd_buffer_io_out_ready = h2m_cmd_buffer_ready_io_ready; // @[Top.scala 185:73]
  assign h2m_cmd_buffer_ready_clock = mmcm_io_CLKOUT1;
  assign h2m_cmd_buffer_ready_reset = ~mmcm_io_LOCKED; // @[Top.scala 184:102]
  assign h2m_cmd_buffer_ready_io_valid = h2m_cmd_buffer_io_out_valid; // @[Top.scala 186:65]
  assign h2m_cmd_buffer_ready_io_complete = h2m_complete_dest_out; // @[Top.scala 187:65]
  assign m2h_start_addr_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign m2h_start_addr_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign m2h_start_addr_src_in = {{30'd0}, d2h_cmd_queue_io_cmd_out_bits_m2h_start_addr}; // @[Top.scala 219:73]
  assign m2h_length_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign m2h_length_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign m2h_length_src_in = d2h_cmd_queue_io_cmd_out_bits_m2h_length; // @[Top.scala 220:73]
  assign m2h_start_pulse_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 41:29]
  assign m2h_start_pulse_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 40:29]
  assign m2h_start_pulse_src_pulse = d2h_cmd_queue_io_cmd_out_ready & d2h_cmd_queue_io_cmd_out_valid; // @[Decoupled.scala 40:37]
  assign m2h_complete_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign m2h_complete_src_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 11:28]
  assign m2h_complete_src_in = m2h_io_complete; // @[Top.scala 216:73]
  assign m2h_last_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign m2h_last_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign m2h_last_src_in = d2h_cmd_queue_io_last; // @[Top.scala 233:81]
  assign m2h_read_count_equal_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign m2h_read_count_equal_src_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 11:28]
  assign m2h_read_count_equal_src_in = m2h_io_read_count_equal; // @[Top.scala 236:65]
  assign c2h_status_clock = qdma_io_pcie_clk; // @[Top.scala 63:39 Top.scala 65:41]
  assign c2h_status_reset = ~pcie_rstn; // @[Top.scala 244:111]
  assign c2h_status_io_c2h_start = c2h_status_start_dest_out; // @[Top.scala 247:73]
  assign c2h_status_io_c2h_status_last = qdma_io_c2h_status_last; // @[Top.scala 249:73]
  assign c2h_status_io_c2h_status_cmp = qdma_io_c2h_status_cmp; // @[Top.scala 248:73]
  assign c2h_status_io_c2h_status_valid = qdma_io_c2h_status_valid; // @[Top.scala 250:73]
  assign c2h_status_io_c2h_status_error = qdma_io_c2h_status_error; // @[Top.scala 251:73]
  assign c2h_status_io_c2h_status_drop = qdma_io_c2h_status_drop; // @[Top.scala 252:73]
  assign c2h_status_start_dest_clk = qdma_io_pcie_clk; // @[Top.scala 63:39 Top.scala 65:41]
  assign c2h_status_start_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign c2h_status_start_src_in = d2h_cmd_queue_io_cmd_out_ready & d2h_cmd_queue_io_cmd_out_valid; // @[Decoupled.scala 40:37]
  assign last_count_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign last_count_src_clk = qdma_io_pcie_clk; // @[Top.scala 63:39 Top.scala 65:41]
  assign last_count_src_in = c2h_status_io_c2h_status_last_count; // @[Top.scala 258:73]
  assign cmp_count_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign cmp_count_src_clk = qdma_io_pcie_clk; // @[Top.scala 63:39 Top.scala 65:41]
  assign cmp_count_src_in = c2h_status_io_c2h_status_cmp_count; // @[Top.scala 260:81]
  assign valid_count_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign valid_count_src_clk = qdma_io_pcie_clk; // @[Top.scala 63:39 Top.scala 65:41]
  assign valid_count_src_in = c2h_status_io_c2h_status_valid_count; // @[Top.scala 262:73]
  assign error_count_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign error_count_src_clk = qdma_io_pcie_clk; // @[Top.scala 63:39 Top.scala 65:41]
  assign error_count_src_in = c2h_status_io_c2h_status_error_count; // @[Top.scala 264:73]
  assign drop_count_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 12:28]
  assign drop_count_src_clk = qdma_io_pcie_clk; // @[Top.scala 63:39 Top.scala 65:41]
  assign drop_count_src_in = c2h_status_io_c2h_status_drop_count; // @[Top.scala 266:73]
  assign h2m_queue_din = qdma_io_h2c_data_bits_data; // @[Top.scala 283:81]
  assign h2m_queue_injectdbiterr = 1'h0;
  assign h2m_queue_injectsbiterr = 1'h0;
  assign h2m_queue_rd_clk = hbmDriver_io_hbm_clk; // @[Top.scala 286:81]
  assign h2m_queue_rd_en = h2m_io_fifo_rden & hbmDriver_io_axi_hbm_0_w_ready; // @[Top.scala 287:87]
  assign h2m_queue_rst = 1'h0; // @[Top.scala 280:81]
  assign h2m_queue_sleep = 1'h0;
  assign h2m_queue_wr_clk = mmcm_io_CLKOUT1; // @[Top.scala 281:81]
  assign h2m_queue_wr_en = qdma_io_h2c_data_valid; // @[Top.scala 282:81]
  assign m2h_queue__din = hbmDriver_io_axi_hbm_0_r_bits_data; // @[Top.scala 299:81]
  assign m2h_queue__injectdbiterr = 1'h0;
  assign m2h_queue__injectsbiterr = 1'h0;
  assign m2h_queue__rd_clk = mmcm_io_CLKOUT1; // @[Top.scala 302:81]
  assign m2h_queue__rd_en = qdma_io_c2h_data_ready & _c2h_io_c2h_cmd_ready_T; // @[Top.scala 303:107]
  assign m2h_queue__rst = 1'h0; // @[Top.scala 296:81]
  assign m2h_queue__sleep = 1'h0;
  assign m2h_queue__wr_clk = hbmDriver_io_hbm_clk; // @[Top.scala 297:73]
  assign m2h_queue__wr_en = hbmDriver_io_axi_hbm_0_r_valid; // @[Top.scala 298:81]
  assign h2m_valid_tmpreg_clock = hbmDriver_io_hbm_clk;
  assign h2m_valid_tmpreg_reset = ~hbm_rstn; // @[Top.scala 289:101]
  assign h2m_valid_tmpreg_io_ready = h2m_io_fifo_rden & hbmDriver_io_axi_hbm_0_w_ready; // @[Top.scala 290:79]
  assign h2m_valid_tmpreg_io_valid = h2m_queue_data_valid; // @[Top.scala 291:73]
  assign m2h_valid_tmpreg_clock = mmcm_io_CLKOUT1;
  assign m2h_valid_tmpreg_reset = ~mmcm_io_LOCKED; // @[Top.scala 305:102]
  assign m2h_valid_tmpreg_io_ready = qdma_io_c2h_data_ready & _c2h_io_c2h_cmd_ready_T; // @[Top.scala 306:99]
  assign m2h_valid_tmpreg_io_valid = m2h_queue__data_valid; // @[Top.scala 307:73]
  assign m2h_queue_empty_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign m2h_queue_empty_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign m2h_queue_empty_src_in = m2h_queue__empty; // @[Top.scala 312:73]
  assign m2h_valid_tmpreg_tom2h_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign m2h_valid_tmpreg_tom2h_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign m2h_valid_tmpreg_tom2h_src_in = m2h_valid_tmpreg_io_tmpreg; // @[Top.scala 315:65]
  assign axicc_s_axi_awaddr = qdma_io_axib_aw_bits_addr; // @[Top.scala 362:57]
  assign axicc_s_axi_awlen = qdma_io_axib_aw_bits_len; // @[Top.scala 363:57]
  assign axicc_s_axi_awsize = qdma_io_axib_aw_bits_size; // @[Top.scala 364:57]
  assign axicc_s_axi_awburst = qdma_io_axib_aw_bits_burst; // @[Top.scala 365:57]
  assign axicc_s_axi_awlock = 1'h0; // @[Top.scala 393:49]
  assign axicc_s_axi_awcache = 4'h0; // @[Top.scala 394:49]
  assign axicc_s_axi_awprot = 3'h0; // @[Top.scala 392:49]
  assign axicc_s_axi_awregion = 4'h0; // @[Top.scala 395:49]
  assign axicc_s_axi_awqos = 4'h0; // @[Top.scala 396:49]
  assign axicc_s_axi_awvalid = qdma_io_axib_aw_valid; // @[Top.scala 366:57]
  assign axicc_s_axi_wdata = qdma_io_axib_w_bits_data; // @[Top.scala 368:57]
  assign axicc_s_axi_wstrb = qdma_io_axib_w_bits_strb; // @[Top.scala 369:57]
  assign axicc_s_axi_wlast = qdma_io_axib_w_bits_last; // @[Top.scala 370:57]
  assign axicc_s_axi_wvalid = qdma_io_axib_w_valid; // @[Top.scala 371:57]
  assign axicc_s_axi_bready = 1'h1; // @[Top.scala 402:49]
  assign axicc_s_axi_araddr = qdma_io_axib_ar_bits_addr; // @[Top.scala 373:57]
  assign axicc_s_axi_arlen = qdma_io_axib_ar_bits_len; // @[Top.scala 374:57]
  assign axicc_s_axi_arsize = qdma_io_axib_ar_bits_size; // @[Top.scala 375:57]
  assign axicc_s_axi_arburst = qdma_io_axib_ar_bits_burst; // @[Top.scala 376:57]
  assign axicc_s_axi_arlock = 1'h0; // @[Top.scala 398:49]
  assign axicc_s_axi_arcache = 4'h0; // @[Top.scala 399:49]
  assign axicc_s_axi_arprot = 3'h0; // @[Top.scala 397:49]
  assign axicc_s_axi_arregion = 4'h0; // @[Top.scala 400:49]
  assign axicc_s_axi_arqos = 4'h0; // @[Top.scala 401:49]
  assign axicc_s_axi_arvalid = qdma_io_axib_ar_valid; // @[Top.scala 377:57]
  assign axicc_s_axi_rready = qdma_io_axib_r_ready; // @[Top.scala 382:57]
  assign axicc_s_axi_aclk = qdma_io_pcie_clk; // @[Top.scala 63:39 Top.scala 65:41]
  assign axicc_s_axi_aresetn = qdma_io_pcie_arstn; // @[Top.scala 64:39 Top.scala 66:41]
  assign axicc_m_axi_aclk = hbmDriver_io_hbm_clk; // @[Top.scala 406:57]
  assign axicc_m_axi_aresetn = hbm_rstn; // @[Top.scala 407:49]
  assign axicc_m_axi_awready = axidwc_s_axi_awready; // @[Top.scala 416:41]
  assign axicc_m_axi_wready = axidwc_s_axi_wready; // @[Top.scala 421:41]
  assign axicc_m_axi_bresp = 2'h0;
  assign axicc_m_axi_bvalid = axidwc_s_axi_bvalid; // @[Top.scala 432:49]
  assign axicc_m_axi_arready = axidwc_s_axi_arready; // @[Top.scala 427:41]
  assign axicc_m_axi_rdata = axidwc_s_axi_rdata; // @[Top.scala 428:41]
  assign axicc_m_axi_rresp = 2'h0;
  assign axicc_m_axi_rlast = axidwc_s_axi_rlast; // @[Top.scala 429:41]
  assign axicc_m_axi_rvalid = axidwc_s_axi_rvalid; // @[Top.scala 430:41]
  assign axidwc_s_axi_awaddr = axicc_m_axi_awaddr[33:0]; // @[Top.scala 411:41]
  assign axidwc_s_axi_awlen = axicc_m_axi_awlen; // @[Top.scala 412:41]
  assign axidwc_s_axi_awsize = axicc_m_axi_awsize; // @[Top.scala 413:41]
  assign axidwc_s_axi_awburst = axicc_m_axi_awburst; // @[Top.scala 414:41]
  assign axidwc_s_axi_awlock = 1'h0; // @[Top.scala 436:49]
  assign axidwc_s_axi_awcache = 4'h0; // @[Top.scala 437:49]
  assign axidwc_s_axi_awprot = 3'h0; // @[Top.scala 435:49]
  assign axidwc_s_axi_awregion = 4'h0; // @[Top.scala 438:49]
  assign axidwc_s_axi_awqos = 4'h0; // @[Top.scala 439:49]
  assign axidwc_s_axi_awvalid = axicc_m_axi_awvalid; // @[Top.scala 415:41]
  assign axidwc_s_axi_wdata = axicc_m_axi_wdata; // @[Top.scala 417:41]
  assign axidwc_s_axi_wstrb = axicc_m_axi_wstrb; // @[Top.scala 418:41]
  assign axidwc_s_axi_wlast = axicc_m_axi_wlast; // @[Top.scala 419:41]
  assign axidwc_s_axi_wvalid = axicc_m_axi_wvalid; // @[Top.scala 420:41]
  assign axidwc_s_axi_bready = 1'h1; // @[Top.scala 445:49]
  assign axidwc_s_axi_araddr = axicc_m_axi_araddr[33:0]; // @[Top.scala 422:41]
  assign axidwc_s_axi_arlen = axicc_m_axi_arlen; // @[Top.scala 423:41]
  assign axidwc_s_axi_arsize = axicc_m_axi_arsize; // @[Top.scala 424:41]
  assign axidwc_s_axi_arburst = axicc_m_axi_arburst; // @[Top.scala 425:41]
  assign axidwc_s_axi_arlock = 1'h0; // @[Top.scala 441:49]
  assign axidwc_s_axi_arcache = 4'h0; // @[Top.scala 442:49]
  assign axidwc_s_axi_arprot = 3'h0; // @[Top.scala 440:49]
  assign axidwc_s_axi_arregion = 4'h0; // @[Top.scala 443:49]
  assign axidwc_s_axi_arqos = 4'h0; // @[Top.scala 444:49]
  assign axidwc_s_axi_arvalid = axicc_m_axi_arvalid; // @[Top.scala 426:41]
  assign axidwc_s_axi_rready = axicc_m_axi_rready; // @[Top.scala 431:41]
  assign axidwc_s_axi_aclk = hbmDriver_io_hbm_clk; // @[Top.scala 408:49]
  assign axidwc_s_axi_aresetn = hbm_rstn; // @[Top.scala 409:49]
  assign axidwc_m_axi_awready = hbmDriver_io_axi_hbm_1_aw_ready; // @[Top.scala 452:41]
  assign axidwc_m_axi_wready = hbmDriver_io_axi_hbm_1_w_ready; // @[Top.scala 457:41]
  assign axidwc_m_axi_bresp = 2'h0;
  assign axidwc_m_axi_bvalid = hbmDriver_io_axi_hbm_1_b_valid; // @[Top.scala 468:49]
  assign axidwc_m_axi_arready = hbmDriver_io_axi_hbm_1_ar_ready; // @[Top.scala 463:41]
  assign axidwc_m_axi_rdata = hbmDriver_io_axi_hbm_1_r_bits_data; // @[Top.scala 464:41]
  assign axidwc_m_axi_rresp = 2'h0;
  assign axidwc_m_axi_rlast = hbmDriver_io_axi_hbm_1_r_bits_last; // @[Top.scala 465:41]
  assign axidwc_m_axi_rvalid = hbmDriver_io_axi_hbm_1_r_valid; // @[Top.scala 466:41]
  assign p2p_counter_clock = hbmDriver_io_hbm_clk;
  assign p2p_counter_reset = ~hbm_rstn; // @[Top.scala 472:85]
  assign p2p_counter_io_start = p2p_counter_io_start_REG; // @[Top.scala 485:49]
  assign p2p_counter_io_length = p2p_length_dest_out; // @[Top.scala 489:49]
  assign p2p_counter_io_wready = hbmDriver_io_axi_hbm_1_w_ready; // @[Top.scala 474:49]
  assign p2p_counter_io_wvalid = hbmDriver_io_axi_hbm_1_w_valid; // @[Top.scala 475:49]
  assign p2p_counter_io_wdatasample = hbmDriver_io_axi_hbm_1_w_bits_data[31:0]; // @[Top.scala 476:87]
  assign p2p_counter_io_p2p_cpt_complete = p2p_cpt_complete_dest_pulse; // @[Top.scala 494:41]
  assign p2p_cpt_addr_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign p2p_cpt_addr_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign p2p_cpt_addr_src_in = {qdma_io_reg_control_92,qdma_io_reg_control_93}; // @[Cat.scala 30:58]
  assign p2p_length_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign p2p_length_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign p2p_length_src_in = qdma_io_reg_control_94; // @[Top.scala 488:49]
  assign p2p_start_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 12:28]
  assign p2p_start_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 11:28]
  assign p2p_start_src_in = p2p_start_io_src_in_REG_2; // @[Top.scala 484:49]
  assign p2p_complete_dest_clk = mmcm_io_CLKOUT1; // @[CDC.scala 41:29]
  assign p2p_complete_src_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 40:29]
  assign p2p_complete_src_pulse = p2p_counter_io_p2p_complete; // @[Top.scala 490:49]
  assign p2p_cpt_complete_dest_clk = hbmDriver_io_hbm_clk; // @[CDC.scala 41:29]
  assign p2p_cpt_complete_src_clk = mmcm_io_CLKOUT1; // @[CDC.scala 40:29]
  assign p2p_cpt_complete_src_pulse = c2h_cpt_io_p2p_cpt_complete; // @[Top.scala 493:41]
  always @(posedge hbmDriver_io_hbm_clk) begin
    hbm_rstn <= hbmDriver_io_hbm_rstn; // @[Top.scala 45:93]
    h2m_io_start_REG <= h2m_start_pulse_dest_pulse; // @[Top.scala 206:128]
    m2h_io_start_REG <= m2h_start_pulse_dest_pulse; // @[Top.scala 224:128]
    p2p_counter_io_start_REG <= p2p_start_dest_out; // @[Top.scala 485:96]
  end
  always @(posedge mmcm_io_CLKOUT1) begin
    h2d_cmd_queue_io_cmd_in_valid_REG <= qdma_io_reg_control_59 == 32'h1; // @[Top.scala 95:157]
    h2d_cmd_queue_io_cmd_in_valid_REG_1 <= h2d_cmd_queue_io_cmd_in_valid_REG; // @[Top.scala 95:133]
    h2d_cmd_queue_io_cmd_in_valid_REG_2 <= h2d_cmd_queue_io_cmd_in_valid_REG_1; // @[Top.scala 95:125]
    h2d_cmd_queue_io_cmd_in_valid_REG_3 <= h2d_cmd_queue_io_cmd_in_valid_REG_2; // @[Top.scala 37:48]
    d2h_cmd_queue_io_cmd_in_valid_REG <= qdma_io_reg_control_79 == 32'h1; // @[Top.scala 120:157]
    d2h_cmd_queue_io_cmd_in_valid_REG_1 <= d2h_cmd_queue_io_cmd_in_valid_REG; // @[Top.scala 120:133]
    d2h_cmd_queue_io_cmd_in_valid_REG_2 <= d2h_cmd_queue_io_cmd_in_valid_REG_1; // @[Top.scala 120:125]
    d2h_cmd_queue_io_cmd_in_valid_REG_3 <= d2h_cmd_queue_io_cmd_in_valid_REG_2; // @[Top.scala 37:48]
    c2h_cpt_io_h2c_start_REG <= h2d_cmd_queue_io_last; // @[Top.scala 37:48]
    c2h_cpt_io_c2h_start_REG <= d2h_cmd_queue_io_last; // @[Top.scala 37:48]
    d2h_cmd_queue_io_h2m_complete_start_REG <= h2d_cmd_queue_io_h2m_complete; // @[Top.scala 37:48]
    if (_T) begin // @[Top.scala 189:121]
      h2m_start_addr_reg <= 34'h0; // @[Top.scala 189:121]
    end else if (_T_9) begin // @[Top.scala 192:43]
      h2m_start_addr_reg <= h2m_cmd_buffer_io_out_bits[65:32]; // @[Top.scala 194:41]
    end
    if (_T) begin // @[Top.scala 190:129]
      h2m_length_reg <= 34'h0; // @[Top.scala 190:129]
    end else if (_T_9) begin // @[Top.scala 192:43]
      h2m_length_reg <= {{2'd0}, h2m_cmd_buffer_io_out_bits[31:0]}; // @[Top.scala 195:41]
    end
    if (_T) begin // @[Top.scala 191:129]
      h2m_last_reg <= 1'h0; // @[Top.scala 191:129]
    end else if (_T_9) begin // @[Top.scala 192:43]
      h2m_last_reg <= h2m_cmd_buffer_io_out_bits[66]; // @[Top.scala 193:41]
    end
    p2p_start_io_src_in_REG <= qdma_io_reg_control_91 == 32'h1; // @[Top.scala 484:131]
    p2p_start_io_src_in_REG_1 <= p2p_start_io_src_in_REG; // @[Top.scala 484:107]
    p2p_start_io_src_in_REG_2 <= p2p_start_io_src_in_REG_1; // @[Top.scala 484:99]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hbm_rstn = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  h2d_cmd_queue_io_cmd_in_valid_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  h2d_cmd_queue_io_cmd_in_valid_REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  h2d_cmd_queue_io_cmd_in_valid_REG_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  h2d_cmd_queue_io_cmd_in_valid_REG_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  d2h_cmd_queue_io_cmd_in_valid_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  d2h_cmd_queue_io_cmd_in_valid_REG_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  d2h_cmd_queue_io_cmd_in_valid_REG_2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  d2h_cmd_queue_io_cmd_in_valid_REG_3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  c2h_cpt_io_h2c_start_REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  c2h_cpt_io_c2h_start_REG = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  d2h_cmd_queue_io_h2m_complete_start_REG = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  h2m_start_addr_reg = _RAND_12[33:0];
  _RAND_13 = {2{`RANDOM}};
  h2m_length_reg = _RAND_13[33:0];
  _RAND_14 = {1{`RANDOM}};
  h2m_last_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  h2m_io_start_REG = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  m2h_io_start_REG = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  p2p_start_io_src_in_REG = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  p2p_start_io_src_in_REG_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  p2p_start_io_src_in_REG_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  p2p_counter_io_start_REG = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
